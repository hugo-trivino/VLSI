
module cpu32 ( power, clk, pc, mem_s, code, write_en, imm_en, branch_en, 
        next_pc );
  output [7:0] pc;
  output [31:0] mem_s;
  input [15:0] code;
  output [7:0] next_pc;
  input power, clk;
  output write_en, imm_en, branch_en;
  wire   n2169, stop_en, jz_en, jnz_en, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         \mypc/temp_pc1[7] , \mypc/temp_pc1[6] , \mypc/temp_pc1[5] ,
         \mypc/temp_pc1[4] , \mypc/temp_pc1[3] , \mypc/temp_pc1[2] ,
         \mypc/temp_pc1[1] , \mypc/temp_pc1[0] , \mypc/temp_pc0[7] ,
         \mypc/temp_pc0[6] , \mypc/temp_pc0[5] , \mypc/temp_pc0[4] ,
         \mypc/temp_pc0[3] , \mypc/temp_pc0[2] , \mypc/temp_pc0[1] ,
         \mypc/temp_pc0[0] , \mypc/inc_pc[7] , \mypc/inc_pc[6] ,
         \mypc/inc_pc[5] , \mypc/inc_pc[4] , \mypc/inc_pc[3] ,
         \mypc/inc_pc[2] , \mypc/inc_pc[1] , \mypc/inc_pc[0] ,
         \mypc/branch_en , \myctl/n6 , \myctl/n5 , \myctl/n4 , \myalu/s0[31] ,
         \myalu/s0[30] , \myalu/s0[29] , \myalu/s0[28] , \myalu/s0[27] ,
         \myalu/s0[26] , \myalu/s0[25] , \myalu/s0[24] , \myalu/s0[23] ,
         \myalu/s0[22] , \myalu/s0[21] , \myalu/s0[20] , \myalu/s0[19] ,
         \myalu/s0[18] , \myalu/s0[17] , \myalu/s0[16] , \myalu/s0[15] ,
         \myalu/s0[14] , \myalu/s0[13] , \myalu/s0[12] , \myalu/s0[11] ,
         \myalu/s0[10] , \myalu/s0[9] , \myalu/s0[8] , \myalu/s0[7] ,
         \myalu/s0[6] , \myalu/s0[5] , \myalu/s0[4] , \myalu/s0[3] ,
         \myalu/s0[2] , \myalu/s0[1] , \myalu/s0[0] , \myalu/s10[31] ,
         \myalu/s10[30] , \myalu/s10[29] , \myalu/s10[28] , \myalu/s10[27] ,
         \myalu/s10[26] , \myalu/s10[25] , \myalu/s10[24] , \myalu/s10[23] ,
         \myalu/s10[22] , \myalu/s10[21] , \myalu/s10[20] , \myalu/s10[19] ,
         \myalu/s10[18] , \myalu/s10[17] , \myalu/s10[16] , \myalu/s10[15] ,
         \myalu/s10[14] , \myalu/s10[13] , \myalu/s10[12] , \myalu/s10[11] ,
         \myalu/s10[10] , \myalu/s10[9] , \myalu/s10[8] , \myalu/s10[7] ,
         \myalu/s10[6] , \myalu/s10[5] , \myalu/s10[4] , \myalu/s10[3] ,
         \myalu/s10[2] , \myalu/s10[1] , \myalu/s10[0] , \myalu/s00[31] ,
         \myalu/s00[30] , \myalu/s00[29] , \myalu/s00[28] , \myalu/s00[27] ,
         \myalu/s00[26] , \myalu/s00[25] , \myalu/s00[24] , \myalu/s00[23] ,
         \myalu/s00[22] , \myalu/s00[21] , \myalu/s00[20] , \myalu/s00[19] ,
         \myalu/s00[18] , \myalu/s00[17] , \myalu/s00[16] , \myalu/s00[15] ,
         \myalu/s00[14] , \myalu/s00[13] , \myalu/s00[12] , \myalu/s00[11] ,
         \myalu/s00[10] , \myalu/s00[9] , \myalu/s00[8] , \myalu/s00[7] ,
         \myalu/s00[6] , \myalu/s00[5] , \myalu/s00[4] , \myalu/s00[3] ,
         \myalu/s00[2] , \myalu/s00[1] , \myalu/s00[0] , \myalu/sxnor[31] ,
         \myalu/sxnor[30] , \myalu/sxnor[29] , \myalu/sxnor[28] ,
         \myalu/sxnor[27] , \myalu/sxnor[26] , \myalu/sxnor[25] ,
         \myalu/sxnor[24] , \myalu/sxnor[23] , \myalu/sxnor[22] ,
         \myalu/sxnor[21] , \myalu/sxnor[20] , \myalu/sxnor[19] ,
         \myalu/sxnor[18] , \myalu/sxnor[17] , \myalu/sxnor[16] ,
         \myalu/sxnor[15] , \myalu/sxnor[14] , \myalu/sxnor[13] ,
         \myalu/sxnor[12] , \myalu/sxnor[11] , \myalu/sxnor[10] ,
         \myalu/sxnor[9] , \myalu/sxnor[8] , \myalu/sxnor[7] ,
         \myalu/sxnor[6] , \myalu/sxnor[5] , \myalu/sxnor[4] ,
         \myalu/sxnor[3] , \myalu/sxnor[2] , \myalu/sxnor[1] ,
         \myalu/sxnor[0] , \myalu/sand[31] , \myalu/sand[30] ,
         \myalu/sand[29] , \myalu/sand[28] , \myalu/sand[27] ,
         \myalu/sand[26] , \myalu/sand[25] , \myalu/sand[24] ,
         \myalu/sand[23] , \myalu/sand[22] , \myalu/sand[21] ,
         \myalu/sand[20] , \myalu/sand[19] , \myalu/sand[18] ,
         \myalu/sand[17] , \myalu/sand[16] , \myalu/sand[15] ,
         \myalu/sand[14] , \myalu/sand[13] , \myalu/sand[12] ,
         \myalu/sand[11] , \myalu/sand[10] , \myalu/sand[9] , \myalu/sand[8] ,
         \myalu/sand[7] , \myalu/sand[6] , \myalu/sand[5] , \myalu/sand[4] ,
         \myalu/sand[3] , \myalu/sand[2] , \myalu/sand[1] , \myalu/sand[0] ,
         \myalu/saddsub[31] , \myalu/saddsub[30] , \myalu/saddsub[29] ,
         \myalu/saddsub[28] , \myalu/saddsub[27] , \myalu/saddsub[26] ,
         \myalu/saddsub[25] , \myalu/saddsub[24] , \myalu/saddsub[23] ,
         \myalu/saddsub[22] , \myalu/saddsub[21] , \myalu/saddsub[20] ,
         \myalu/saddsub[19] , \myalu/saddsub[18] , \myalu/saddsub[17] ,
         \myalu/saddsub[16] , \myalu/saddsub[15] , \myalu/saddsub[14] ,
         \myalu/saddsub[13] , \myalu/saddsub[12] , \myalu/saddsub[11] ,
         \myalu/saddsub[10] , \myalu/saddsub[9] , \myalu/saddsub[8] ,
         \myalu/saddsub[7] , \myalu/saddsub[6] , \myalu/saddsub[5] ,
         \myalu/saddsub[4] , \myalu/saddsub[3] , \myalu/saddsub[2] ,
         \myalu/saddsub[1] , \myalu/saddsub[0] , \myalu/ssr[31] ,
         \myalu/ssr[30] , \myalu/ssr[29] , \myalu/ssr[28] , \myalu/ssr[27] ,
         \myalu/ssr[26] , \myalu/ssr[25] , \myalu/ssr[24] , \myalu/ssr[23] ,
         \myalu/ssr[22] , \myalu/ssr[21] , \myalu/ssr[20] , \myalu/ssr[19] ,
         \myalu/ssr[18] , \myalu/ssr[17] , \myalu/ssr[16] , \myalu/ssr[15] ,
         \myalu/ssr[14] , \myalu/ssr[13] , \myalu/ssr[12] , \myalu/ssr[11] ,
         \myalu/ssr[10] , \myalu/ssr[9] , \myalu/ssr[8] , \myalu/ssr[7] ,
         \myalu/ssr[6] , \myalu/ssr[5] , \myalu/ssr[4] , \myalu/ssr[3] ,
         \myalu/ssr[2] , \myalu/ssr[1] , \myalu/ssr[0] , \myalu/ssl[31] ,
         \myalu/ssl[30] , \myalu/ssl[29] , \myalu/ssl[28] , \myalu/ssl[27] ,
         \myalu/ssl[26] , \myalu/ssl[25] , \myalu/ssl[24] , \myalu/ssl[23] ,
         \myalu/ssl[22] , \myalu/ssl[21] , \myalu/ssl[20] , \myalu/ssl[19] ,
         \myalu/ssl[18] , \myalu/ssl[17] , \myalu/ssl[16] , \myalu/ssl[15] ,
         \myalu/ssl[14] , \myalu/ssl[13] , \myalu/ssl[12] , \myalu/ssl[11] ,
         \myalu/ssl[10] , \myalu/ssl[9] , \myalu/ssl[8] , \myalu/ssl[7] ,
         \myalu/ssl[6] , \myalu/ssl[5] , \myalu/ssl[4] , \myalu/ssl[3] ,
         \myalu/ssl[2] , \myalu/ssl[1] , \myalu/ssl[0] , \myram/sel_s[15] ,
         \myram/sel_s[14] , \myram/sel_s[13] , \myram/sel_s[12] ,
         \myram/sel_s[11] , \myram/sel_s[10] , \myram/sel_s[9] ,
         \myram/sel_s[8] , \myram/sel_s[7] , \myram/sel_s[6] ,
         \myram/sel_s[5] , \myram/sel_s[4] , \myram/sel_s[3] ,
         \myram/sel_s[2] , \myram/sel_s[1] , \myram/sel_s[0] ,
         \myram/sel_b[15] , \myram/sel_b[14] , \myram/sel_b[13] ,
         \myram/sel_b[12] , \myram/sel_b[11] , \myram/sel_b[10] ,
         \myram/sel_b[9] , \myram/sel_b[8] , \myram/sel_b[7] ,
         \myram/sel_b[6] , \myram/sel_b[5] , \myram/sel_b[4] ,
         \myram/sel_b[3] , \myram/sel_b[2] , \myram/sel_b[1] ,
         \myram/sel_b[0] , \myram/sel_a[15] , \myram/sel_a[14] ,
         \myram/sel_a[13] , \myram/sel_a[12] , \myram/sel_a[11] ,
         \myram/sel_a[10] , \myram/sel_a[9] , \myram/sel_a[8] ,
         \myram/sel_a[7] , \myram/sel_a[6] , \myram/sel_a[5] ,
         \myram/sel_a[4] , \myram/sel_a[3] , \myram/sel_a[2] ,
         \myram/sel_a[1] , \myram/sel_a[0] , \myalu/mysll/s4[0] ,
         \myalu/mysll/s4[1] , \myalu/mysll/s4[2] , \myalu/mysll/s4[3] ,
         \myalu/mysll/s4[4] , \myalu/mysll/s4[5] , \myalu/mysll/s4[6] ,
         \myalu/mysll/s4[7] , \myalu/mysll/s4[8] , \myalu/mysll/s4[9] ,
         \myalu/mysll/s4[10] , \myalu/mysll/s4[11] , \myalu/mysll/s4[12] ,
         \myalu/mysll/s4[13] , \myalu/mysll/s4[14] , \myalu/mysll/s4[15] ,
         \myalu/mysll/s4[16] , \myalu/mysll/s4[17] , \myalu/mysll/s4[18] ,
         \myalu/mysll/s4[19] , \myalu/mysll/s4[20] , \myalu/mysll/s4[21] ,
         \myalu/mysll/s4[22] , \myalu/mysll/s4[23] , \myalu/mysll/s4[24] ,
         \myalu/mysll/s4[25] , \myalu/mysll/s4[26] , \myalu/mysll/s4[27] ,
         \myalu/mysll/s4[28] , \myalu/mysll/s4[29] , \myalu/mysll/s4[30] ,
         \myalu/mysll/s4[31] , \myalu/mysll/s3[0] , \myalu/mysll/s3[1] ,
         \myalu/mysll/s3[2] , \myalu/mysll/s3[3] , \myalu/mysll/s3[4] ,
         \myalu/mysll/s3[5] , \myalu/mysll/s3[6] , \myalu/mysll/s3[7] ,
         \myalu/mysll/s3[8] , \myalu/mysll/s3[9] , \myalu/mysll/s3[10] ,
         \myalu/mysll/s3[11] , \myalu/mysll/s3[12] , \myalu/mysll/s3[13] ,
         \myalu/mysll/s3[14] , \myalu/mysll/s3[15] , \myalu/mysll/s3[16] ,
         \myalu/mysll/s3[17] , \myalu/mysll/s3[18] , \myalu/mysll/s3[19] ,
         \myalu/mysll/s3[20] , \myalu/mysll/s3[21] , \myalu/mysll/s3[22] ,
         \myalu/mysll/s3[23] , \myalu/mysll/s3[24] , \myalu/mysll/s3[25] ,
         \myalu/mysll/s3[26] , \myalu/mysll/s3[27] , \myalu/mysll/s3[28] ,
         \myalu/mysll/s3[29] , \myalu/mysll/s3[30] , \myalu/mysll/s3[31] ,
         \myalu/mysll/s2[0] , \myalu/mysll/s2[1] , \myalu/mysll/s2[2] ,
         \myalu/mysll/s2[3] , \myalu/mysll/s2[4] , \myalu/mysll/s2[5] ,
         \myalu/mysll/s2[6] , \myalu/mysll/s2[7] , \myalu/mysll/s2[8] ,
         \myalu/mysll/s2[9] , \myalu/mysll/s2[10] , \myalu/mysll/s2[11] ,
         \myalu/mysll/s2[12] , \myalu/mysll/s2[13] , \myalu/mysll/s2[14] ,
         \myalu/mysll/s2[15] , \myalu/mysll/s2[16] , \myalu/mysll/s2[17] ,
         \myalu/mysll/s2[18] , \myalu/mysll/s2[19] , \myalu/mysll/s2[20] ,
         \myalu/mysll/s2[21] , \myalu/mysll/s2[22] , \myalu/mysll/s2[23] ,
         \myalu/mysll/s2[24] , \myalu/mysll/s2[25] , \myalu/mysll/s2[26] ,
         \myalu/mysll/s2[27] , \myalu/mysll/s2[28] , \myalu/mysll/s2[29] ,
         \myalu/mysll/s2[30] , \myalu/mysll/s2[31] , \myalu/mysll/s1[0] ,
         \myalu/mysll/s1[1] , \myalu/mysll/s1[2] , \myalu/mysll/s1[3] ,
         \myalu/mysll/s1[4] , \myalu/mysll/s1[5] , \myalu/mysll/s1[6] ,
         \myalu/mysll/s1[7] , \myalu/mysll/s1[8] , \myalu/mysll/s1[9] ,
         \myalu/mysll/s1[10] , \myalu/mysll/s1[11] , \myalu/mysll/s1[12] ,
         \myalu/mysll/s1[13] , \myalu/mysll/s1[14] , \myalu/mysll/s1[15] ,
         \myalu/mysll/s1[16] , \myalu/mysll/s1[17] , \myalu/mysll/s1[18] ,
         \myalu/mysll/s1[19] , \myalu/mysll/s1[20] , \myalu/mysll/s1[21] ,
         \myalu/mysll/s1[22] , \myalu/mysll/s1[23] , \myalu/mysll/s1[24] ,
         \myalu/mysll/s1[25] , \myalu/mysll/s1[26] , \myalu/mysll/s1[27] ,
         \myalu/mysll/s1[28] , \myalu/mysll/s1[29] , \myalu/mysll/s1[30] ,
         \myalu/mysll/s1[31] , \myalu/mysrl/s4[0] , \myalu/mysrl/s4[1] ,
         \myalu/mysrl/s4[2] , \myalu/mysrl/s4[3] , \myalu/mysrl/s4[4] ,
         \myalu/mysrl/s4[5] , \myalu/mysrl/s4[6] , \myalu/mysrl/s4[7] ,
         \myalu/mysrl/s4[8] , \myalu/mysrl/s4[9] , \myalu/mysrl/s4[10] ,
         \myalu/mysrl/s4[11] , \myalu/mysrl/s4[12] , \myalu/mysrl/s4[13] ,
         \myalu/mysrl/s4[14] , \myalu/mysrl/s4[15] , \myalu/mysrl/s4[16] ,
         \myalu/mysrl/s4[17] , \myalu/mysrl/s4[18] , \myalu/mysrl/s4[19] ,
         \myalu/mysrl/s4[20] , \myalu/mysrl/s4[21] , \myalu/mysrl/s4[22] ,
         \myalu/mysrl/s4[23] , \myalu/mysrl/s4[24] , \myalu/mysrl/s4[25] ,
         \myalu/mysrl/s4[26] , \myalu/mysrl/s4[27] , \myalu/mysrl/s4[28] ,
         \myalu/mysrl/s4[29] , \myalu/mysrl/s4[30] , \myalu/mysrl/s4[31] ,
         \myalu/mysrl/s3[0] , \myalu/mysrl/s3[1] , \myalu/mysrl/s3[2] ,
         \myalu/mysrl/s3[3] , \myalu/mysrl/s3[4] , \myalu/mysrl/s3[5] ,
         \myalu/mysrl/s3[6] , \myalu/mysrl/s3[7] , \myalu/mysrl/s3[8] ,
         \myalu/mysrl/s3[9] , \myalu/mysrl/s3[10] , \myalu/mysrl/s3[11] ,
         \myalu/mysrl/s3[12] , \myalu/mysrl/s3[13] , \myalu/mysrl/s3[14] ,
         \myalu/mysrl/s3[15] , \myalu/mysrl/s3[16] , \myalu/mysrl/s3[17] ,
         \myalu/mysrl/s3[18] , \myalu/mysrl/s3[19] , \myalu/mysrl/s3[20] ,
         \myalu/mysrl/s3[21] , \myalu/mysrl/s3[22] , \myalu/mysrl/s3[23] ,
         \myalu/mysrl/s3[24] , \myalu/mysrl/s3[25] , \myalu/mysrl/s3[26] ,
         \myalu/mysrl/s3[27] , \myalu/mysrl/s3[28] , \myalu/mysrl/s3[29] ,
         \myalu/mysrl/s3[30] , \myalu/mysrl/s3[31] , \myalu/mysrl/s2[0] ,
         \myalu/mysrl/s2[1] , \myalu/mysrl/s2[2] , \myalu/mysrl/s2[3] ,
         \myalu/mysrl/s2[4] , \myalu/mysrl/s2[5] , \myalu/mysrl/s2[6] ,
         \myalu/mysrl/s2[7] , \myalu/mysrl/s2[8] , \myalu/mysrl/s2[9] ,
         \myalu/mysrl/s2[10] , \myalu/mysrl/s2[11] , \myalu/mysrl/s2[12] ,
         \myalu/mysrl/s2[13] , \myalu/mysrl/s2[14] , \myalu/mysrl/s2[15] ,
         \myalu/mysrl/s2[16] , \myalu/mysrl/s2[17] , \myalu/mysrl/s2[18] ,
         \myalu/mysrl/s2[19] , \myalu/mysrl/s2[20] , \myalu/mysrl/s2[21] ,
         \myalu/mysrl/s2[22] , \myalu/mysrl/s2[23] , \myalu/mysrl/s2[24] ,
         \myalu/mysrl/s2[25] , \myalu/mysrl/s2[26] , \myalu/mysrl/s2[27] ,
         \myalu/mysrl/s2[28] , \myalu/mysrl/s2[29] , \myalu/mysrl/s2[30] ,
         \myalu/mysrl/s2[31] , \myalu/mysrl/s1[0] , \myalu/mysrl/s1[1] ,
         \myalu/mysrl/s1[2] , \myalu/mysrl/s1[3] , \myalu/mysrl/s1[4] ,
         \myalu/mysrl/s1[5] , \myalu/mysrl/s1[6] , \myalu/mysrl/s1[7] ,
         \myalu/mysrl/s1[8] , \myalu/mysrl/s1[9] , \myalu/mysrl/s1[10] ,
         \myalu/mysrl/s1[11] , \myalu/mysrl/s1[12] , \myalu/mysrl/s1[13] ,
         \myalu/mysrl/s1[14] , \myalu/mysrl/s1[15] , \myalu/mysrl/s1[16] ,
         \myalu/mysrl/s1[17] , \myalu/mysrl/s1[18] , \myalu/mysrl/s1[19] ,
         \myalu/mysrl/s1[20] , \myalu/mysrl/s1[21] , \myalu/mysrl/s1[22] ,
         \myalu/mysrl/s1[23] , \myalu/mysrl/s1[24] , \myalu/mysrl/s1[25] ,
         \myalu/mysrl/s1[26] , \myalu/mysrl/s1[27] , \myalu/mysrl/s1[28] ,
         \myalu/mysrl/s1[29] , \myalu/mysrl/s1[30] , \myalu/mysrl/s1[31] ,
         \myalu/myadder/xb[31] , \myalu/myadder/xb[30] ,
         \myalu/myadder/xb[29] , \myalu/myadder/xb[28] ,
         \myalu/myadder/xb[27] , \myalu/myadder/xb[26] ,
         \myalu/myadder/xb[25] , \myalu/myadder/xb[24] ,
         \myalu/myadder/xb[23] , \myalu/myadder/xb[22] ,
         \myalu/myadder/xb[21] , \myalu/myadder/xb[20] ,
         \myalu/myadder/xb[19] , \myalu/myadder/xb[18] ,
         \myalu/myadder/xb[17] , \myalu/myadder/xb[16] ,
         \myalu/myadder/xb[15] , \myalu/myadder/xb[14] ,
         \myalu/myadder/xb[13] , \myalu/myadder/xb[12] ,
         \myalu/myadder/xb[11] , \myalu/myadder/xb[10] , \myalu/myadder/xb[9] ,
         \myalu/myadder/xb[8] , \myalu/myadder/xb[7] , \myalu/myadder/xb[6] ,
         \myalu/myadder/xb[5] , \myalu/myadder/xb[4] , \myalu/myadder/xb[3] ,
         \myalu/myadder/xb[2] , \myalu/myadder/xb[1] , \myalu/myadder/xb[0] ,
         \myram/da/en1 , \myram/da/en0 , \myram/m0/mux_out[31] ,
         \myram/m0/mux_out[30] , \myram/m0/mux_out[29] ,
         \myram/m0/mux_out[28] , \myram/m0/mux_out[27] ,
         \myram/m0/mux_out[26] , \myram/m0/mux_out[25] ,
         \myram/m0/mux_out[24] , \myram/m0/mux_out[23] ,
         \myram/m0/mux_out[22] , \myram/m0/mux_out[21] ,
         \myram/m0/mux_out[20] , \myram/m0/mux_out[19] ,
         \myram/m0/mux_out[18] , \myram/m0/mux_out[17] ,
         \myram/m0/mux_out[16] , \myram/m0/mux_out[15] ,
         \myram/m0/mux_out[14] , \myram/m0/mux_out[13] ,
         \myram/m0/mux_out[12] , \myram/m0/mux_out[11] ,
         \myram/m0/mux_out[10] , \myram/m0/mux_out[9] , \myram/m0/mux_out[8] ,
         \myram/m0/mux_out[7] , \myram/m0/mux_out[6] , \myram/m0/mux_out[5] ,
         \myram/m0/mux_out[4] , \myram/m0/mux_out[3] , \myram/m0/mux_out[2] ,
         \myram/m0/mux_out[1] , \myram/m0/mux_out[0] , \myram/m0/dout[0] ,
         \myram/m0/dout[1] , \myram/m0/dout[2] , \myram/m0/dout[3] ,
         \myram/m0/dout[4] , \myram/m0/dout[5] , \myram/m0/dout[6] ,
         \myram/m0/dout[7] , \myram/m0/dout[8] , \myram/m0/dout[9] ,
         \myram/m0/dout[10] , \myram/m0/dout[11] , \myram/m0/dout[12] ,
         \myram/m0/dout[13] , \myram/m0/dout[14] , \myram/m0/dout[15] ,
         \myram/m0/dout[16] , \myram/m0/dout[17] , \myram/m0/dout[18] ,
         \myram/m0/dout[19] , \myram/m0/dout[20] , \myram/m0/dout[21] ,
         \myram/m0/dout[22] , \myram/m0/dout[23] , \myram/m0/dout[24] ,
         \myram/m0/dout[25] , \myram/m0/dout[26] , \myram/m0/dout[27] ,
         \myram/m0/dout[28] , \myram/m0/dout[29] , \myram/m0/dout[30] ,
         \myram/m0/dout[31] , \myram/m1/mux_out[31] , \myram/m1/mux_out[30] ,
         \myram/m1/mux_out[29] , \myram/m1/mux_out[28] ,
         \myram/m1/mux_out[27] , \myram/m1/mux_out[26] ,
         \myram/m1/mux_out[25] , \myram/m1/mux_out[24] ,
         \myram/m1/mux_out[23] , \myram/m1/mux_out[22] ,
         \myram/m1/mux_out[21] , \myram/m1/mux_out[20] ,
         \myram/m1/mux_out[19] , \myram/m1/mux_out[18] ,
         \myram/m1/mux_out[17] , \myram/m1/mux_out[16] ,
         \myram/m1/mux_out[15] , \myram/m1/mux_out[14] ,
         \myram/m1/mux_out[13] , \myram/m1/mux_out[12] ,
         \myram/m1/mux_out[11] , \myram/m1/mux_out[10] , \myram/m1/mux_out[9] ,
         \myram/m1/mux_out[8] , \myram/m1/mux_out[7] , \myram/m1/mux_out[6] ,
         \myram/m1/mux_out[5] , \myram/m1/mux_out[4] , \myram/m1/mux_out[3] ,
         \myram/m1/mux_out[2] , \myram/m1/mux_out[1] , \myram/m1/mux_out[0] ,
         \myram/m1/dout[0] , \myram/m1/dout[1] , \myram/m1/dout[2] ,
         \myram/m1/dout[3] , \myram/m1/dout[4] , \myram/m1/dout[5] ,
         \myram/m1/dout[6] , \myram/m1/dout[7] , \myram/m1/dout[8] ,
         \myram/m1/dout[9] , \myram/m1/dout[10] , \myram/m1/dout[11] ,
         \myram/m1/dout[12] , \myram/m1/dout[13] , \myram/m1/dout[14] ,
         \myram/m1/dout[15] , \myram/m1/dout[16] , \myram/m1/dout[17] ,
         \myram/m1/dout[18] , \myram/m1/dout[19] , \myram/m1/dout[20] ,
         \myram/m1/dout[21] , \myram/m1/dout[22] , \myram/m1/dout[23] ,
         \myram/m1/dout[24] , \myram/m1/dout[25] , \myram/m1/dout[26] ,
         \myram/m1/dout[27] , \myram/m1/dout[28] , \myram/m1/dout[29] ,
         \myram/m1/dout[30] , \myram/m1/dout[31] , \alu_out/m0/n3 ,
         \myalu/myadder/myadder/c31 , \myalu/myadder/myadder/c30 ,
         \myalu/myadder/myadder/c29 , \myalu/myadder/myadder/c28 ,
         \myalu/myadder/myadder/c27 , \myalu/myadder/myadder/c26 ,
         \myalu/myadder/myadder/c25 , \myalu/myadder/myadder/c24 ,
         \myalu/myadder/myadder/c23 , \myalu/myadder/myadder/c22 ,
         \myalu/myadder/myadder/c21 , \myalu/myadder/myadder/c20 ,
         \myalu/myadder/myadder/c19 , \myalu/myadder/myadder/c18 ,
         \myalu/myadder/myadder/c17 , \myalu/myadder/myadder/c16 ,
         \myalu/myadder/myadder/c15 , \myalu/myadder/myadder/c14 ,
         \myalu/myadder/myadder/c13 , \myalu/myadder/myadder/c12 ,
         \myalu/myadder/myadder/c11 , \myalu/myadder/myadder/c10 ,
         \myalu/myadder/myadder/c9 , \myalu/myadder/myadder/c8 ,
         \myalu/myadder/myadder/c7 , \myalu/myadder/myadder/c6 ,
         \myalu/myadder/myadder/c5 , \myalu/myadder/myadder/c4 ,
         \myalu/myadder/myadder/c3 , \myalu/myadder/myadder/c2 ,
         \myalu/myadder/myadder/c1 , \myram/da/d0/en1 , \myram/ds/en1 ,
         \myram/ds/en0 , \myram/db/en1 , \myram/m15/mux_out[31] ,
         \myram/m15/mux_out[30] , \myram/m15/mux_out[29] ,
         \myram/m15/mux_out[28] , \myram/m15/mux_out[27] ,
         \myram/m15/mux_out[26] , \myram/m15/mux_out[25] ,
         \myram/m15/mux_out[24] , \myram/m15/mux_out[23] ,
         \myram/m15/mux_out[22] , \myram/m15/mux_out[21] ,
         \myram/m15/mux_out[20] , \myram/m15/mux_out[19] ,
         \myram/m15/mux_out[18] , \myram/m15/mux_out[17] ,
         \myram/m15/mux_out[16] , \myram/m15/mux_out[15] ,
         \myram/m15/mux_out[14] , \myram/m15/mux_out[13] ,
         \myram/m15/mux_out[12] , \myram/m15/mux_out[11] ,
         \myram/m15/mux_out[10] , \myram/m15/mux_out[9] ,
         \myram/m15/mux_out[8] , \myram/m15/mux_out[7] ,
         \myram/m15/mux_out[6] , \myram/m15/mux_out[5] ,
         \myram/m15/mux_out[4] , \myram/m15/mux_out[3] ,
         \myram/m15/mux_out[2] , \myram/m15/mux_out[1] ,
         \myram/m15/mux_out[0] , \myram/m15/dout[0] , \myram/m15/dout[1] ,
         \myram/m15/dout[2] , \myram/m15/dout[3] , \myram/m15/dout[4] ,
         \myram/m15/dout[5] , \myram/m15/dout[6] , \myram/m15/dout[7] ,
         \myram/m15/dout[8] , \myram/m15/dout[9] , \myram/m15/dout[10] ,
         \myram/m15/dout[11] , \myram/m15/dout[12] , \myram/m15/dout[13] ,
         \myram/m15/dout[14] , \myram/m15/dout[15] , \myram/m15/dout[16] ,
         \myram/m15/dout[17] , \myram/m15/dout[18] , \myram/m15/dout[19] ,
         \myram/m15/dout[20] , \myram/m15/dout[21] , \myram/m15/dout[22] ,
         \myram/m15/dout[23] , \myram/m15/dout[24] , \myram/m15/dout[25] ,
         \myram/m15/dout[26] , \myram/m15/dout[27] , \myram/m15/dout[28] ,
         \myram/m15/dout[29] , \myram/m15/dout[30] , \myram/m15/dout[31] ,
         \myram/m14/mux_out[31] , \myram/m14/mux_out[30] ,
         \myram/m14/mux_out[29] , \myram/m14/mux_out[28] ,
         \myram/m14/mux_out[27] , \myram/m14/mux_out[26] ,
         \myram/m14/mux_out[25] , \myram/m14/mux_out[24] ,
         \myram/m14/mux_out[23] , \myram/m14/mux_out[22] ,
         \myram/m14/mux_out[21] , \myram/m14/mux_out[20] ,
         \myram/m14/mux_out[19] , \myram/m14/mux_out[18] ,
         \myram/m14/mux_out[17] , \myram/m14/mux_out[16] ,
         \myram/m14/mux_out[15] , \myram/m14/mux_out[14] ,
         \myram/m14/mux_out[13] , \myram/m14/mux_out[12] ,
         \myram/m14/mux_out[11] , \myram/m14/mux_out[10] ,
         \myram/m14/mux_out[9] , \myram/m14/mux_out[8] ,
         \myram/m14/mux_out[7] , \myram/m14/mux_out[6] ,
         \myram/m14/mux_out[5] , \myram/m14/mux_out[4] ,
         \myram/m14/mux_out[3] , \myram/m14/mux_out[2] ,
         \myram/m14/mux_out[1] , \myram/m14/mux_out[0] , \myram/m14/dout[0] ,
         \myram/m14/dout[1] , \myram/m14/dout[2] , \myram/m14/dout[3] ,
         \myram/m14/dout[4] , \myram/m14/dout[5] , \myram/m14/dout[6] ,
         \myram/m14/dout[7] , \myram/m14/dout[8] , \myram/m14/dout[9] ,
         \myram/m14/dout[10] , \myram/m14/dout[11] , \myram/m14/dout[12] ,
         \myram/m14/dout[13] , \myram/m14/dout[14] , \myram/m14/dout[15] ,
         \myram/m14/dout[16] , \myram/m14/dout[17] , \myram/m14/dout[18] ,
         \myram/m14/dout[19] , \myram/m14/dout[20] , \myram/m14/dout[21] ,
         \myram/m14/dout[22] , \myram/m14/dout[23] , \myram/m14/dout[24] ,
         \myram/m14/dout[25] , \myram/m14/dout[26] , \myram/m14/dout[27] ,
         \myram/m14/dout[28] , \myram/m14/dout[29] , \myram/m14/dout[30] ,
         \myram/m14/dout[31] , \myram/m13/mux_out[31] ,
         \myram/m13/mux_out[30] , \myram/m13/mux_out[29] ,
         \myram/m13/mux_out[28] , \myram/m13/mux_out[27] ,
         \myram/m13/mux_out[26] , \myram/m13/mux_out[25] ,
         \myram/m13/mux_out[24] , \myram/m13/mux_out[23] ,
         \myram/m13/mux_out[22] , \myram/m13/mux_out[21] ,
         \myram/m13/mux_out[20] , \myram/m13/mux_out[19] ,
         \myram/m13/mux_out[18] , \myram/m13/mux_out[17] ,
         \myram/m13/mux_out[16] , \myram/m13/mux_out[15] ,
         \myram/m13/mux_out[14] , \myram/m13/mux_out[13] ,
         \myram/m13/mux_out[12] , \myram/m13/mux_out[11] ,
         \myram/m13/mux_out[10] , \myram/m13/mux_out[9] ,
         \myram/m13/mux_out[8] , \myram/m13/mux_out[7] ,
         \myram/m13/mux_out[6] , \myram/m13/mux_out[5] ,
         \myram/m13/mux_out[4] , \myram/m13/mux_out[3] ,
         \myram/m13/mux_out[2] , \myram/m13/mux_out[1] ,
         \myram/m13/mux_out[0] , \myram/m13/dout[0] , \myram/m13/dout[1] ,
         \myram/m13/dout[2] , \myram/m13/dout[3] , \myram/m13/dout[4] ,
         \myram/m13/dout[5] , \myram/m13/dout[6] , \myram/m13/dout[7] ,
         \myram/m13/dout[8] , \myram/m13/dout[9] , \myram/m13/dout[10] ,
         \myram/m13/dout[11] , \myram/m13/dout[12] , \myram/m13/dout[13] ,
         \myram/m13/dout[14] , \myram/m13/dout[15] , \myram/m13/dout[16] ,
         \myram/m13/dout[17] , \myram/m13/dout[18] , \myram/m13/dout[19] ,
         \myram/m13/dout[20] , \myram/m13/dout[21] , \myram/m13/dout[22] ,
         \myram/m13/dout[23] , \myram/m13/dout[24] , \myram/m13/dout[25] ,
         \myram/m13/dout[26] , \myram/m13/dout[27] , \myram/m13/dout[28] ,
         \myram/m13/dout[29] , \myram/m13/dout[30] , \myram/m13/dout[31] ,
         \myram/m12/mux_out[31] , \myram/m12/mux_out[30] ,
         \myram/m12/mux_out[29] , \myram/m12/mux_out[28] ,
         \myram/m12/mux_out[27] , \myram/m12/mux_out[26] ,
         \myram/m12/mux_out[25] , \myram/m12/mux_out[24] ,
         \myram/m12/mux_out[23] , \myram/m12/mux_out[22] ,
         \myram/m12/mux_out[21] , \myram/m12/mux_out[20] ,
         \myram/m12/mux_out[19] , \myram/m12/mux_out[18] ,
         \myram/m12/mux_out[17] , \myram/m12/mux_out[16] ,
         \myram/m12/mux_out[15] , \myram/m12/mux_out[14] ,
         \myram/m12/mux_out[13] , \myram/m12/mux_out[12] ,
         \myram/m12/mux_out[11] , \myram/m12/mux_out[10] ,
         \myram/m12/mux_out[9] , \myram/m12/mux_out[8] ,
         \myram/m12/mux_out[7] , \myram/m12/mux_out[6] ,
         \myram/m12/mux_out[5] , \myram/m12/mux_out[4] ,
         \myram/m12/mux_out[3] , \myram/m12/mux_out[2] ,
         \myram/m12/mux_out[1] , \myram/m12/mux_out[0] , \myram/m12/dout[0] ,
         \myram/m12/dout[1] , \myram/m12/dout[2] , \myram/m12/dout[3] ,
         \myram/m12/dout[4] , \myram/m12/dout[5] , \myram/m12/dout[6] ,
         \myram/m12/dout[7] , \myram/m12/dout[8] , \myram/m12/dout[9] ,
         \myram/m12/dout[10] , \myram/m12/dout[11] , \myram/m12/dout[12] ,
         \myram/m12/dout[13] , \myram/m12/dout[14] , \myram/m12/dout[15] ,
         \myram/m12/dout[16] , \myram/m12/dout[17] , \myram/m12/dout[18] ,
         \myram/m12/dout[19] , \myram/m12/dout[20] , \myram/m12/dout[21] ,
         \myram/m12/dout[22] , \myram/m12/dout[23] , \myram/m12/dout[24] ,
         \myram/m12/dout[25] , \myram/m12/dout[26] , \myram/m12/dout[27] ,
         \myram/m12/dout[28] , \myram/m12/dout[29] , \myram/m12/dout[30] ,
         \myram/m12/dout[31] , \myram/m11/mux_out[31] ,
         \myram/m11/mux_out[30] , \myram/m11/mux_out[29] ,
         \myram/m11/mux_out[28] , \myram/m11/mux_out[27] ,
         \myram/m11/mux_out[26] , \myram/m11/mux_out[25] ,
         \myram/m11/mux_out[24] , \myram/m11/mux_out[23] ,
         \myram/m11/mux_out[22] , \myram/m11/mux_out[21] ,
         \myram/m11/mux_out[20] , \myram/m11/mux_out[19] ,
         \myram/m11/mux_out[18] , \myram/m11/mux_out[17] ,
         \myram/m11/mux_out[16] , \myram/m11/mux_out[15] ,
         \myram/m11/mux_out[14] , \myram/m11/mux_out[13] ,
         \myram/m11/mux_out[12] , \myram/m11/mux_out[11] ,
         \myram/m11/mux_out[10] , \myram/m11/mux_out[9] ,
         \myram/m11/mux_out[8] , \myram/m11/mux_out[7] ,
         \myram/m11/mux_out[6] , \myram/m11/mux_out[5] ,
         \myram/m11/mux_out[4] , \myram/m11/mux_out[3] ,
         \myram/m11/mux_out[2] , \myram/m11/mux_out[1] ,
         \myram/m11/mux_out[0] , \myram/m11/dout[0] , \myram/m11/dout[1] ,
         \myram/m11/dout[2] , \myram/m11/dout[3] , \myram/m11/dout[4] ,
         \myram/m11/dout[5] , \myram/m11/dout[6] , \myram/m11/dout[7] ,
         \myram/m11/dout[8] , \myram/m11/dout[9] , \myram/m11/dout[10] ,
         \myram/m11/dout[11] , \myram/m11/dout[12] , \myram/m11/dout[13] ,
         \myram/m11/dout[14] , \myram/m11/dout[15] , \myram/m11/dout[16] ,
         \myram/m11/dout[17] , \myram/m11/dout[18] , \myram/m11/dout[19] ,
         \myram/m11/dout[20] , \myram/m11/dout[21] , \myram/m11/dout[22] ,
         \myram/m11/dout[23] , \myram/m11/dout[24] , \myram/m11/dout[25] ,
         \myram/m11/dout[26] , \myram/m11/dout[27] , \myram/m11/dout[28] ,
         \myram/m11/dout[29] , \myram/m11/dout[30] , \myram/m11/dout[31] ,
         \myram/m10/mux_out[31] , \myram/m10/mux_out[30] ,
         \myram/m10/mux_out[29] , \myram/m10/mux_out[28] ,
         \myram/m10/mux_out[27] , \myram/m10/mux_out[26] ,
         \myram/m10/mux_out[25] , \myram/m10/mux_out[24] ,
         \myram/m10/mux_out[23] , \myram/m10/mux_out[22] ,
         \myram/m10/mux_out[21] , \myram/m10/mux_out[20] ,
         \myram/m10/mux_out[19] , \myram/m10/mux_out[18] ,
         \myram/m10/mux_out[17] , \myram/m10/mux_out[16] ,
         \myram/m10/mux_out[15] , \myram/m10/mux_out[14] ,
         \myram/m10/mux_out[13] , \myram/m10/mux_out[12] ,
         \myram/m10/mux_out[11] , \myram/m10/mux_out[10] ,
         \myram/m10/mux_out[9] , \myram/m10/mux_out[8] ,
         \myram/m10/mux_out[7] , \myram/m10/mux_out[6] ,
         \myram/m10/mux_out[5] , \myram/m10/mux_out[4] ,
         \myram/m10/mux_out[3] , \myram/m10/mux_out[2] ,
         \myram/m10/mux_out[1] , \myram/m10/mux_out[0] , \myram/m10/dout[0] ,
         \myram/m10/dout[1] , \myram/m10/dout[2] , \myram/m10/dout[3] ,
         \myram/m10/dout[4] , \myram/m10/dout[5] , \myram/m10/dout[6] ,
         \myram/m10/dout[7] , \myram/m10/dout[8] , \myram/m10/dout[9] ,
         \myram/m10/dout[10] , \myram/m10/dout[11] , \myram/m10/dout[12] ,
         \myram/m10/dout[13] , \myram/m10/dout[14] , \myram/m10/dout[15] ,
         \myram/m10/dout[16] , \myram/m10/dout[17] , \myram/m10/dout[18] ,
         \myram/m10/dout[19] , \myram/m10/dout[20] , \myram/m10/dout[21] ,
         \myram/m10/dout[22] , \myram/m10/dout[23] , \myram/m10/dout[24] ,
         \myram/m10/dout[25] , \myram/m10/dout[26] , \myram/m10/dout[27] ,
         \myram/m10/dout[28] , \myram/m10/dout[29] , \myram/m10/dout[30] ,
         \myram/m10/dout[31] , \myram/m9/mux_out[31] , \myram/m9/mux_out[30] ,
         \myram/m9/mux_out[29] , \myram/m9/mux_out[28] ,
         \myram/m9/mux_out[27] , \myram/m9/mux_out[26] ,
         \myram/m9/mux_out[25] , \myram/m9/mux_out[24] ,
         \myram/m9/mux_out[23] , \myram/m9/mux_out[22] ,
         \myram/m9/mux_out[21] , \myram/m9/mux_out[20] ,
         \myram/m9/mux_out[19] , \myram/m9/mux_out[18] ,
         \myram/m9/mux_out[17] , \myram/m9/mux_out[16] ,
         \myram/m9/mux_out[15] , \myram/m9/mux_out[14] ,
         \myram/m9/mux_out[13] , \myram/m9/mux_out[12] ,
         \myram/m9/mux_out[11] , \myram/m9/mux_out[10] , \myram/m9/mux_out[9] ,
         \myram/m9/mux_out[8] , \myram/m9/mux_out[7] , \myram/m9/mux_out[6] ,
         \myram/m9/mux_out[5] , \myram/m9/mux_out[4] , \myram/m9/mux_out[3] ,
         \myram/m9/mux_out[2] , \myram/m9/mux_out[1] , \myram/m9/mux_out[0] ,
         \myram/m9/dout[0] , \myram/m9/dout[1] , \myram/m9/dout[2] ,
         \myram/m9/dout[3] , \myram/m9/dout[4] , \myram/m9/dout[5] ,
         \myram/m9/dout[6] , \myram/m9/dout[7] , \myram/m9/dout[8] ,
         \myram/m9/dout[9] , \myram/m9/dout[10] , \myram/m9/dout[11] ,
         \myram/m9/dout[12] , \myram/m9/dout[13] , \myram/m9/dout[14] ,
         \myram/m9/dout[15] , \myram/m9/dout[16] , \myram/m9/dout[17] ,
         \myram/m9/dout[18] , \myram/m9/dout[19] , \myram/m9/dout[20] ,
         \myram/m9/dout[21] , \myram/m9/dout[22] , \myram/m9/dout[23] ,
         \myram/m9/dout[24] , \myram/m9/dout[25] , \myram/m9/dout[26] ,
         \myram/m9/dout[27] , \myram/m9/dout[28] , \myram/m9/dout[29] ,
         \myram/m9/dout[30] , \myram/m9/dout[31] , \myram/m8/mux_out[31] ,
         \myram/m8/mux_out[30] , \myram/m8/mux_out[29] ,
         \myram/m8/mux_out[28] , \myram/m8/mux_out[27] ,
         \myram/m8/mux_out[26] , \myram/m8/mux_out[25] ,
         \myram/m8/mux_out[24] , \myram/m8/mux_out[23] ,
         \myram/m8/mux_out[22] , \myram/m8/mux_out[21] ,
         \myram/m8/mux_out[20] , \myram/m8/mux_out[19] ,
         \myram/m8/mux_out[18] , \myram/m8/mux_out[17] ,
         \myram/m8/mux_out[16] , \myram/m8/mux_out[15] ,
         \myram/m8/mux_out[14] , \myram/m8/mux_out[13] ,
         \myram/m8/mux_out[12] , \myram/m8/mux_out[11] ,
         \myram/m8/mux_out[10] , \myram/m8/mux_out[9] , \myram/m8/mux_out[8] ,
         \myram/m8/mux_out[7] , \myram/m8/mux_out[6] , \myram/m8/mux_out[5] ,
         \myram/m8/mux_out[4] , \myram/m8/mux_out[3] , \myram/m8/mux_out[2] ,
         \myram/m8/mux_out[1] , \myram/m8/mux_out[0] , \myram/m8/dout[0] ,
         \myram/m8/dout[1] , \myram/m8/dout[2] , \myram/m8/dout[3] ,
         \myram/m8/dout[4] , \myram/m8/dout[5] , \myram/m8/dout[6] ,
         \myram/m8/dout[7] , \myram/m8/dout[8] , \myram/m8/dout[9] ,
         \myram/m8/dout[10] , \myram/m8/dout[11] , \myram/m8/dout[12] ,
         \myram/m8/dout[13] , \myram/m8/dout[14] , \myram/m8/dout[15] ,
         \myram/m8/dout[16] , \myram/m8/dout[17] , \myram/m8/dout[18] ,
         \myram/m8/dout[19] , \myram/m8/dout[20] , \myram/m8/dout[21] ,
         \myram/m8/dout[22] , \myram/m8/dout[23] , \myram/m8/dout[24] ,
         \myram/m8/dout[25] , \myram/m8/dout[26] , \myram/m8/dout[27] ,
         \myram/m8/dout[28] , \myram/m8/dout[29] , \myram/m8/dout[30] ,
         \myram/m8/dout[31] , \myram/m7/mux_out[31] , \myram/m7/mux_out[30] ,
         \myram/m7/mux_out[29] , \myram/m7/mux_out[28] ,
         \myram/m7/mux_out[27] , \myram/m7/mux_out[26] ,
         \myram/m7/mux_out[25] , \myram/m7/mux_out[24] ,
         \myram/m7/mux_out[23] , \myram/m7/mux_out[22] ,
         \myram/m7/mux_out[21] , \myram/m7/mux_out[20] ,
         \myram/m7/mux_out[19] , \myram/m7/mux_out[18] ,
         \myram/m7/mux_out[17] , \myram/m7/mux_out[16] ,
         \myram/m7/mux_out[15] , \myram/m7/mux_out[14] ,
         \myram/m7/mux_out[13] , \myram/m7/mux_out[12] ,
         \myram/m7/mux_out[11] , \myram/m7/mux_out[10] , \myram/m7/mux_out[9] ,
         \myram/m7/mux_out[8] , \myram/m7/mux_out[7] , \myram/m7/mux_out[6] ,
         \myram/m7/mux_out[5] , \myram/m7/mux_out[4] , \myram/m7/mux_out[3] ,
         \myram/m7/mux_out[2] , \myram/m7/mux_out[1] , \myram/m7/mux_out[0] ,
         \myram/m7/dout[0] , \myram/m7/dout[1] , \myram/m7/dout[2] ,
         \myram/m7/dout[3] , \myram/m7/dout[4] , \myram/m7/dout[5] ,
         \myram/m7/dout[6] , \myram/m7/dout[7] , \myram/m7/dout[8] ,
         \myram/m7/dout[9] , \myram/m7/dout[10] , \myram/m7/dout[11] ,
         \myram/m7/dout[12] , \myram/m7/dout[13] , \myram/m7/dout[14] ,
         \myram/m7/dout[15] , \myram/m7/dout[16] , \myram/m7/dout[17] ,
         \myram/m7/dout[18] , \myram/m7/dout[19] , \myram/m7/dout[20] ,
         \myram/m7/dout[21] , \myram/m7/dout[22] , \myram/m7/dout[23] ,
         \myram/m7/dout[24] , \myram/m7/dout[25] , \myram/m7/dout[26] ,
         \myram/m7/dout[27] , \myram/m7/dout[28] , \myram/m7/dout[29] ,
         \myram/m7/dout[30] , \myram/m7/dout[31] , \myram/m6/mux_out[31] ,
         \myram/m6/mux_out[30] , \myram/m6/mux_out[29] ,
         \myram/m6/mux_out[28] , \myram/m6/mux_out[27] ,
         \myram/m6/mux_out[26] , \myram/m6/mux_out[25] ,
         \myram/m6/mux_out[24] , \myram/m6/mux_out[23] ,
         \myram/m6/mux_out[22] , \myram/m6/mux_out[21] ,
         \myram/m6/mux_out[20] , \myram/m6/mux_out[19] ,
         \myram/m6/mux_out[18] , \myram/m6/mux_out[17] ,
         \myram/m6/mux_out[16] , \myram/m6/mux_out[15] ,
         \myram/m6/mux_out[14] , \myram/m6/mux_out[13] ,
         \myram/m6/mux_out[12] , \myram/m6/mux_out[11] ,
         \myram/m6/mux_out[10] , \myram/m6/mux_out[9] , \myram/m6/mux_out[8] ,
         \myram/m6/mux_out[7] , \myram/m6/mux_out[6] , \myram/m6/mux_out[5] ,
         \myram/m6/mux_out[4] , \myram/m6/mux_out[3] , \myram/m6/mux_out[2] ,
         \myram/m6/mux_out[1] , \myram/m6/mux_out[0] , \myram/m6/dout[0] ,
         \myram/m6/dout[1] , \myram/m6/dout[2] , \myram/m6/dout[3] ,
         \myram/m6/dout[4] , \myram/m6/dout[5] , \myram/m6/dout[6] ,
         \myram/m6/dout[7] , \myram/m6/dout[8] , \myram/m6/dout[9] ,
         \myram/m6/dout[10] , \myram/m6/dout[11] , \myram/m6/dout[12] ,
         \myram/m6/dout[13] , \myram/m6/dout[14] , \myram/m6/dout[15] ,
         \myram/m6/dout[16] , \myram/m6/dout[17] , \myram/m6/dout[18] ,
         \myram/m6/dout[19] , \myram/m6/dout[20] , \myram/m6/dout[21] ,
         \myram/m6/dout[22] , \myram/m6/dout[23] , \myram/m6/dout[24] ,
         \myram/m6/dout[25] , \myram/m6/dout[26] , \myram/m6/dout[27] ,
         \myram/m6/dout[28] , \myram/m6/dout[29] , \myram/m6/dout[30] ,
         \myram/m6/dout[31] , \myram/m5/mux_out[31] , \myram/m5/mux_out[30] ,
         \myram/m5/mux_out[29] , \myram/m5/mux_out[28] ,
         \myram/m5/mux_out[27] , \myram/m5/mux_out[26] ,
         \myram/m5/mux_out[25] , \myram/m5/mux_out[24] ,
         \myram/m5/mux_out[23] , \myram/m5/mux_out[22] ,
         \myram/m5/mux_out[21] , \myram/m5/mux_out[20] ,
         \myram/m5/mux_out[19] , \myram/m5/mux_out[18] ,
         \myram/m5/mux_out[17] , \myram/m5/mux_out[16] ,
         \myram/m5/mux_out[15] , \myram/m5/mux_out[14] ,
         \myram/m5/mux_out[13] , \myram/m5/mux_out[12] ,
         \myram/m5/mux_out[11] , \myram/m5/mux_out[10] , \myram/m5/mux_out[9] ,
         \myram/m5/mux_out[8] , \myram/m5/mux_out[7] , \myram/m5/mux_out[6] ,
         \myram/m5/mux_out[5] , \myram/m5/mux_out[4] , \myram/m5/mux_out[3] ,
         \myram/m5/mux_out[2] , \myram/m5/mux_out[1] , \myram/m5/mux_out[0] ,
         \myram/m5/dout[0] , \myram/m5/dout[1] , \myram/m5/dout[2] ,
         \myram/m5/dout[3] , \myram/m5/dout[4] , \myram/m5/dout[5] ,
         \myram/m5/dout[6] , \myram/m5/dout[7] , \myram/m5/dout[8] ,
         \myram/m5/dout[9] , \myram/m5/dout[10] , \myram/m5/dout[11] ,
         \myram/m5/dout[12] , \myram/m5/dout[13] , \myram/m5/dout[14] ,
         \myram/m5/dout[15] , \myram/m5/dout[16] , \myram/m5/dout[17] ,
         \myram/m5/dout[18] , \myram/m5/dout[19] , \myram/m5/dout[20] ,
         \myram/m5/dout[21] , \myram/m5/dout[22] , \myram/m5/dout[23] ,
         \myram/m5/dout[24] , \myram/m5/dout[25] , \myram/m5/dout[26] ,
         \myram/m5/dout[27] , \myram/m5/dout[28] , \myram/m5/dout[29] ,
         \myram/m5/dout[30] , \myram/m5/dout[31] , \myram/m4/mux_out[31] ,
         \myram/m4/mux_out[30] , \myram/m4/mux_out[29] ,
         \myram/m4/mux_out[28] , \myram/m4/mux_out[27] ,
         \myram/m4/mux_out[26] , \myram/m4/mux_out[25] ,
         \myram/m4/mux_out[24] , \myram/m4/mux_out[23] ,
         \myram/m4/mux_out[22] , \myram/m4/mux_out[21] ,
         \myram/m4/mux_out[20] , \myram/m4/mux_out[19] ,
         \myram/m4/mux_out[18] , \myram/m4/mux_out[17] ,
         \myram/m4/mux_out[16] , \myram/m4/mux_out[15] ,
         \myram/m4/mux_out[14] , \myram/m4/mux_out[13] ,
         \myram/m4/mux_out[12] , \myram/m4/mux_out[11] ,
         \myram/m4/mux_out[10] , \myram/m4/mux_out[9] , \myram/m4/mux_out[8] ,
         \myram/m4/mux_out[7] , \myram/m4/mux_out[6] , \myram/m4/mux_out[5] ,
         \myram/m4/mux_out[4] , \myram/m4/mux_out[3] , \myram/m4/mux_out[2] ,
         \myram/m4/mux_out[1] , \myram/m4/mux_out[0] , \myram/m4/dout[0] ,
         \myram/m4/dout[1] , \myram/m4/dout[2] , \myram/m4/dout[3] ,
         \myram/m4/dout[4] , \myram/m4/dout[5] , \myram/m4/dout[6] ,
         \myram/m4/dout[7] , \myram/m4/dout[8] , \myram/m4/dout[9] ,
         \myram/m4/dout[10] , \myram/m4/dout[11] , \myram/m4/dout[12] ,
         \myram/m4/dout[13] , \myram/m4/dout[14] , \myram/m4/dout[15] ,
         \myram/m4/dout[16] , \myram/m4/dout[17] , \myram/m4/dout[18] ,
         \myram/m4/dout[19] , \myram/m4/dout[20] , \myram/m4/dout[21] ,
         \myram/m4/dout[22] , \myram/m4/dout[23] , \myram/m4/dout[24] ,
         \myram/m4/dout[25] , \myram/m4/dout[26] , \myram/m4/dout[27] ,
         \myram/m4/dout[28] , \myram/m4/dout[29] , \myram/m4/dout[30] ,
         \myram/m4/dout[31] , \myram/m3/mux_out[31] , \myram/m3/mux_out[30] ,
         \myram/m3/mux_out[29] , \myram/m3/mux_out[28] ,
         \myram/m3/mux_out[27] , \myram/m3/mux_out[26] ,
         \myram/m3/mux_out[25] , \myram/m3/mux_out[24] ,
         \myram/m3/mux_out[23] , \myram/m3/mux_out[22] ,
         \myram/m3/mux_out[21] , \myram/m3/mux_out[20] ,
         \myram/m3/mux_out[19] , \myram/m3/mux_out[18] ,
         \myram/m3/mux_out[17] , \myram/m3/mux_out[16] ,
         \myram/m3/mux_out[15] , \myram/m3/mux_out[14] ,
         \myram/m3/mux_out[13] , \myram/m3/mux_out[12] ,
         \myram/m3/mux_out[11] , \myram/m3/mux_out[10] , \myram/m3/mux_out[9] ,
         \myram/m3/mux_out[8] , \myram/m3/mux_out[7] , \myram/m3/mux_out[6] ,
         \myram/m3/mux_out[5] , \myram/m3/mux_out[4] , \myram/m3/mux_out[3] ,
         \myram/m3/mux_out[2] , \myram/m3/mux_out[1] , \myram/m3/mux_out[0] ,
         \myram/m3/dout[0] , \myram/m3/dout[1] , \myram/m3/dout[2] ,
         \myram/m3/dout[3] , \myram/m3/dout[4] , \myram/m3/dout[5] ,
         \myram/m3/dout[6] , \myram/m3/dout[7] , \myram/m3/dout[8] ,
         \myram/m3/dout[9] , \myram/m3/dout[10] , \myram/m3/dout[11] ,
         \myram/m3/dout[12] , \myram/m3/dout[13] , \myram/m3/dout[14] ,
         \myram/m3/dout[15] , \myram/m3/dout[16] , \myram/m3/dout[17] ,
         \myram/m3/dout[18] , \myram/m3/dout[19] , \myram/m3/dout[20] ,
         \myram/m3/dout[21] , \myram/m3/dout[22] , \myram/m3/dout[23] ,
         \myram/m3/dout[24] , \myram/m3/dout[25] , \myram/m3/dout[26] ,
         \myram/m3/dout[27] , \myram/m3/dout[28] , \myram/m3/dout[29] ,
         \myram/m3/dout[30] , \myram/m3/dout[31] , \myram/m2/mux_out[31] ,
         \myram/m2/mux_out[30] , \myram/m2/mux_out[29] ,
         \myram/m2/mux_out[28] , \myram/m2/mux_out[27] ,
         \myram/m2/mux_out[26] , \myram/m2/mux_out[25] ,
         \myram/m2/mux_out[24] , \myram/m2/mux_out[23] ,
         \myram/m2/mux_out[22] , \myram/m2/mux_out[21] ,
         \myram/m2/mux_out[20] , \myram/m2/mux_out[19] ,
         \myram/m2/mux_out[18] , \myram/m2/mux_out[17] ,
         \myram/m2/mux_out[16] , \myram/m2/mux_out[15] ,
         \myram/m2/mux_out[14] , \myram/m2/mux_out[13] ,
         \myram/m2/mux_out[12] , \myram/m2/mux_out[11] ,
         \myram/m2/mux_out[10] , \myram/m2/mux_out[9] , \myram/m2/mux_out[8] ,
         \myram/m2/mux_out[7] , \myram/m2/mux_out[6] , \myram/m2/mux_out[5] ,
         \myram/m2/mux_out[4] , \myram/m2/mux_out[3] , \myram/m2/mux_out[2] ,
         \myram/m2/mux_out[1] , \myram/m2/mux_out[0] , \myram/m2/dout[0] ,
         \myram/m2/dout[1] , \myram/m2/dout[2] , \myram/m2/dout[3] ,
         \myram/m2/dout[4] , \myram/m2/dout[5] , \myram/m2/dout[6] ,
         \myram/m2/dout[7] , \myram/m2/dout[8] , \myram/m2/dout[9] ,
         \myram/m2/dout[10] , \myram/m2/dout[11] , \myram/m2/dout[12] ,
         \myram/m2/dout[13] , \myram/m2/dout[14] , \myram/m2/dout[15] ,
         \myram/m2/dout[16] , \myram/m2/dout[17] , \myram/m2/dout[18] ,
         \myram/m2/dout[19] , \myram/m2/dout[20] , \myram/m2/dout[21] ,
         \myram/m2/dout[22] , \myram/m2/dout[23] , \myram/m2/dout[24] ,
         \myram/m2/dout[25] , \myram/m2/dout[26] , \myram/m2/dout[27] ,
         \myram/m2/dout[28] , \myram/m2/dout[29] , \myram/m2/dout[30] ,
         \myram/m2/dout[31] , \myram/ds/d1/en1 , \myram/ds/d0/en1 ,
         \myram/db/d1/en1 , \myram/db/d0/en1 , \myram/da/d1/en1 , n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n125, n126, n128, n129, n132, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168;
  wire   [3:0] addr_s;
  wire   [3:0] addr_a;
  wire   [3:0] addr_b;
  wire   [2:0] alu_op;
  wire   [31:0] alu_s;
  tri   [31:0] a;
  tri   [31:0] b;
  assign addr_s[3] = code[11];
  assign addr_s[2] = code[10];
  assign addr_s[1] = code[9];
  assign addr_s[0] = code[8];
  assign addr_a[2] = code[6];
  assign addr_a[1] = code[5];
  assign addr_a[0] = code[4];
  assign addr_b[2] = code[2];
  assign addr_b[1] = code[1];
  assign addr_b[0] = code[0];
  assign alu_op[2] = code[14];
  assign alu_op[1] = code[13];
  assign alu_op[0] = code[12];
  assign branch_en = \mypc/branch_en ;
  assign \myram/da/en1  = code[7];
  assign \myram/db/en1  = code[3];

  AOI22X1 U15 ( .A(jz_en), .B(n2), .C(jnz_en), .D(n4), .Y(n3) );
  NAND3X1 U16 ( .A(n7), .B(n8), .C(n9), .Y(n6) );
  NOR3X1 U17 ( .A(n12), .B(a[21]), .C(a[20]), .Y(n11) );
  NOR3X1 U18 ( .A(n13), .B(a[18]), .C(a[17]), .Y(n10) );
  NOR3X1 U19 ( .A(n14), .B(a[14]), .C(a[13]), .Y(n8) );
  NOR3X1 U20 ( .A(n15), .B(a[10]), .C(a[0]), .Y(n7) );
  NAND3X1 U21 ( .A(n16), .B(n17), .C(n18), .Y(n5) );
  NOR3X1 U22 ( .A(n21), .B(a[7]), .C(a[6]), .Y(n20) );
  NOR3X1 U23 ( .A(n22), .B(a[3]), .C(a[31]), .Y(n19) );
  NOR3X1 U24 ( .A(n23), .B(a[29]), .C(a[28]), .Y(n17) );
  NOR3X1 U25 ( .A(n24), .B(a[25]), .C(a[24]), .Y(n16) );
  NOR3X1 \myctl/U10  ( .A(n126), .B(n310), .C(n313), .Y(imm_en) );
  NOR3X1 \myctl/U9  ( .A(n126), .B(alu_op[1]), .C(n312), .Y(jnz_en) );
  NOR3X1 \myctl/U8  ( .A(n126), .B(alu_op[1]), .C(n310), .Y(jz_en) );
  NOR3X1 \myctl/U6  ( .A(n61), .B(n312), .C(n314), .Y(stop_en) );
  NAND3X1 \myctl/U5  ( .A(n312), .B(n314), .C(alu_op[1]), .Y(\myctl/n4 ) );
  XOR2X1 \myalu/myadder/U32  ( .A(n310), .B(b[0]), .Y(\myalu/myadder/xb[0] )
         );
  XOR2X1 \myalu/myadder/U31  ( .A(n310), .B(b[10]), .Y(\myalu/myadder/xb[10] )
         );
  XOR2X1 \myalu/myadder/U30  ( .A(n310), .B(b[11]), .Y(\myalu/myadder/xb[11] )
         );
  XOR2X1 \myalu/myadder/U29  ( .A(n310), .B(b[12]), .Y(\myalu/myadder/xb[12] )
         );
  XOR2X1 \myalu/myadder/U28  ( .A(n310), .B(b[13]), .Y(\myalu/myadder/xb[13] )
         );
  XOR2X1 \myalu/myadder/U27  ( .A(n310), .B(b[14]), .Y(\myalu/myadder/xb[14] )
         );
  XOR2X1 \myalu/myadder/U26  ( .A(n309), .B(b[15]), .Y(\myalu/myadder/xb[15] )
         );
  XOR2X1 \myalu/myadder/U25  ( .A(n309), .B(b[16]), .Y(\myalu/myadder/xb[16] )
         );
  XOR2X1 \myalu/myadder/U24  ( .A(n309), .B(b[17]), .Y(\myalu/myadder/xb[17] )
         );
  XOR2X1 \myalu/myadder/U23  ( .A(n309), .B(b[18]), .Y(\myalu/myadder/xb[18] )
         );
  XOR2X1 \myalu/myadder/U22  ( .A(n309), .B(b[19]), .Y(\myalu/myadder/xb[19] )
         );
  XOR2X1 \myalu/myadder/U21  ( .A(n309), .B(n62), .Y(\myalu/myadder/xb[1] ) );
  XOR2X1 \myalu/myadder/U20  ( .A(n309), .B(b[20]), .Y(\myalu/myadder/xb[20] )
         );
  XOR2X1 \myalu/myadder/U19  ( .A(n309), .B(b[21]), .Y(\myalu/myadder/xb[21] )
         );
  XOR2X1 \myalu/myadder/U18  ( .A(n309), .B(b[22]), .Y(\myalu/myadder/xb[22] )
         );
  XOR2X1 \myalu/myadder/U17  ( .A(n309), .B(b[23]), .Y(\myalu/myadder/xb[23] )
         );
  XOR2X1 \myalu/myadder/U16  ( .A(n309), .B(b[24]), .Y(\myalu/myadder/xb[24] )
         );
  XOR2X1 \myalu/myadder/U15  ( .A(n309), .B(b[25]), .Y(\myalu/myadder/xb[25] )
         );
  XOR2X1 \myalu/myadder/U14  ( .A(n308), .B(b[26]), .Y(\myalu/myadder/xb[26] )
         );
  XOR2X1 \myalu/myadder/U13  ( .A(n309), .B(b[27]), .Y(\myalu/myadder/xb[27] )
         );
  XOR2X1 \myalu/myadder/U12  ( .A(n308), .B(b[28]), .Y(\myalu/myadder/xb[28] )
         );
  XOR2X1 \myalu/myadder/U11  ( .A(n308), .B(b[29]), .Y(\myalu/myadder/xb[29] )
         );
  XOR2X1 \myalu/myadder/U10  ( .A(n308), .B(n25), .Y(\myalu/myadder/xb[2] ) );
  XOR2X1 \myalu/myadder/U9  ( .A(n308), .B(b[30]), .Y(\myalu/myadder/xb[30] )
         );
  XOR2X1 \myalu/myadder/U8  ( .A(n308), .B(b[31]), .Y(\myalu/myadder/xb[31] )
         );
  XOR2X1 \myalu/myadder/U7  ( .A(n308), .B(b[3]), .Y(\myalu/myadder/xb[3] ) );
  XOR2X1 \myalu/myadder/U6  ( .A(n308), .B(b[4]), .Y(\myalu/myadder/xb[4] ) );
  XOR2X1 \myalu/myadder/U5  ( .A(n308), .B(b[5]), .Y(\myalu/myadder/xb[5] ) );
  XOR2X1 \myalu/myadder/U4  ( .A(n308), .B(b[6]), .Y(\myalu/myadder/xb[6] ) );
  XOR2X1 \myalu/myadder/U3  ( .A(n308), .B(b[7]), .Y(\myalu/myadder/xb[7] ) );
  XOR2X1 \myalu/myadder/U2  ( .A(n308), .B(b[8]), .Y(\myalu/myadder/xb[8] ) );
  XOR2X1 \myalu/myadder/U1  ( .A(n308), .B(b[9]), .Y(\myalu/myadder/xb[9] ) );
  XNOR2X1 \myalu/myxnor/U32  ( .A(n129), .B(a[0]), .Y(\myalu/sxnor[0] ) );
  XNOR2X1 \myalu/myxnor/U31  ( .A(n62), .B(a[1]), .Y(\myalu/sxnor[1] ) );
  XNOR2X1 \myalu/myxnor/U30  ( .A(n25), .B(a[2]), .Y(\myalu/sxnor[2] ) );
  XNOR2X1 \myalu/myxnor/U29  ( .A(b[3]), .B(a[3]), .Y(\myalu/sxnor[3] ) );
  XNOR2X1 \myalu/myxnor/U28  ( .A(b[4]), .B(a[4]), .Y(\myalu/sxnor[4] ) );
  XNOR2X1 \myalu/myxnor/U27  ( .A(b[5]), .B(a[5]), .Y(\myalu/sxnor[5] ) );
  XNOR2X1 \myalu/myxnor/U26  ( .A(b[6]), .B(a[6]), .Y(\myalu/sxnor[6] ) );
  XNOR2X1 \myalu/myxnor/U25  ( .A(b[7]), .B(a[7]), .Y(\myalu/sxnor[7] ) );
  XNOR2X1 \myalu/myxnor/U24  ( .A(b[8]), .B(a[8]), .Y(\myalu/sxnor[8] ) );
  XNOR2X1 \myalu/myxnor/U23  ( .A(b[9]), .B(a[9]), .Y(\myalu/sxnor[9] ) );
  XNOR2X1 \myalu/myxnor/U22  ( .A(b[10]), .B(a[10]), .Y(\myalu/sxnor[10] ) );
  XNOR2X1 \myalu/myxnor/U21  ( .A(b[11]), .B(a[11]), .Y(\myalu/sxnor[11] ) );
  XNOR2X1 \myalu/myxnor/U20  ( .A(b[12]), .B(a[12]), .Y(\myalu/sxnor[12] ) );
  XNOR2X1 \myalu/myxnor/U19  ( .A(b[13]), .B(a[13]), .Y(\myalu/sxnor[13] ) );
  XNOR2X1 \myalu/myxnor/U18  ( .A(b[14]), .B(a[14]), .Y(\myalu/sxnor[14] ) );
  XNOR2X1 \myalu/myxnor/U17  ( .A(b[15]), .B(a[15]), .Y(\myalu/sxnor[15] ) );
  XNOR2X1 \myalu/myxnor/U16  ( .A(b[16]), .B(a[16]), .Y(\myalu/sxnor[16] ) );
  XNOR2X1 \myalu/myxnor/U15  ( .A(b[17]), .B(a[17]), .Y(\myalu/sxnor[17] ) );
  XNOR2X1 \myalu/myxnor/U14  ( .A(b[18]), .B(a[18]), .Y(\myalu/sxnor[18] ) );
  XNOR2X1 \myalu/myxnor/U13  ( .A(b[19]), .B(a[19]), .Y(\myalu/sxnor[19] ) );
  XNOR2X1 \myalu/myxnor/U12  ( .A(b[20]), .B(a[20]), .Y(\myalu/sxnor[20] ) );
  XNOR2X1 \myalu/myxnor/U11  ( .A(b[21]), .B(a[21]), .Y(\myalu/sxnor[21] ) );
  XNOR2X1 \myalu/myxnor/U10  ( .A(b[22]), .B(a[22]), .Y(\myalu/sxnor[22] ) );
  XNOR2X1 \myalu/myxnor/U9  ( .A(b[23]), .B(a[23]), .Y(\myalu/sxnor[23] ) );
  XNOR2X1 \myalu/myxnor/U8  ( .A(b[24]), .B(a[24]), .Y(\myalu/sxnor[24] ) );
  XNOR2X1 \myalu/myxnor/U7  ( .A(b[25]), .B(a[25]), .Y(\myalu/sxnor[25] ) );
  XNOR2X1 \myalu/myxnor/U6  ( .A(b[26]), .B(a[26]), .Y(\myalu/sxnor[26] ) );
  XNOR2X1 \myalu/myxnor/U5  ( .A(b[27]), .B(a[27]), .Y(\myalu/sxnor[27] ) );
  XNOR2X1 \myalu/myxnor/U4  ( .A(b[28]), .B(a[28]), .Y(\myalu/sxnor[28] ) );
  XNOR2X1 \myalu/myxnor/U3  ( .A(b[29]), .B(a[29]), .Y(\myalu/sxnor[29] ) );
  XNOR2X1 \myalu/myxnor/U2  ( .A(b[30]), .B(a[30]), .Y(\myalu/sxnor[30] ) );
  XNOR2X1 \myalu/myxnor/U1  ( .A(b[31]), .B(a[31]), .Y(\myalu/sxnor[31] ) );
  AOI22X1 \alu_out/m0/U3  ( .A(alu_s[0]), .B(n315), .C(imm_en), .D(n205), .Y(
        \alu_out/m0/n3 ) );
  DFFPOSX1 \mypc/d/d0/q_reg  ( .D(next_pc[0]), .CLK(clk), .Q(pc[0]) );
  NOR3X1 \myram/da/d0/d0/U7  ( .A(n192), .B(n208), .C(n207), .Y(
        \myram/sel_a[0] ) );
  NOR3X1 \myram/da/d0/d0/U6  ( .A(n829), .B(n208), .C(n192), .Y(
        \myram/sel_a[1] ) );
  NOR3X1 \myram/da/d0/d0/U5  ( .A(n828), .B(n207), .C(n192), .Y(
        \myram/sel_a[2] ) );
  NOR3X1 \myram/da/d0/d0/U4  ( .A(n828), .B(n192), .C(n829), .Y(
        \myram/sel_a[3] ) );
  TBUFX2 \myram/m0/ta/t0/b1  ( .A(n343), .EN(\myram/sel_a[0] ), .Y(a[0]) );
  AOI22X1 \myram/m15/m0/m31/U3  ( .A(\myram/m15/dout[31] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(n132), .Y(n2168) );
  AOI22X1 \myram/m15/m0/m30/U3  ( .A(\myram/m15/dout[30] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[30]), .Y(n2167) );
  AOI22X1 \myram/m15/m0/m29/U3  ( .A(\myram/m15/dout[29] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[29]), .Y(n2166) );
  AOI22X1 \myram/m15/m0/m28/U3  ( .A(\myram/m15/dout[28] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[28]), .Y(n2165) );
  AOI22X1 \myram/m15/m0/m27/U3  ( .A(\myram/m15/dout[27] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[27]), .Y(n2164) );
  AOI22X1 \myram/m15/m0/m26/U3  ( .A(\myram/m15/dout[26] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[26]), .Y(n2163) );
  AOI22X1 \myram/m15/m0/m25/U3  ( .A(\myram/m15/dout[25] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[25]), .Y(n2162) );
  AOI22X1 \myram/m15/m0/m24/U3  ( .A(\myram/m15/dout[24] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[24]), .Y(n2161) );
  AOI22X1 \myram/m15/m0/m23/U3  ( .A(\myram/m15/dout[23] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[23]), .Y(n2160) );
  AOI22X1 \myram/m15/m0/m22/U3  ( .A(\myram/m15/dout[22] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[22]), .Y(n2159) );
  AOI22X1 \myram/m15/m0/m21/U3  ( .A(\myram/m15/dout[21] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[21]), .Y(n2158) );
  AOI22X1 \myram/m15/m0/m20/U3  ( .A(\myram/m15/dout[20] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[20]), .Y(n2157) );
  AOI22X1 \myram/m15/m0/m19/U3  ( .A(\myram/m15/dout[19] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[19]), .Y(n2156) );
  AOI22X1 \myram/m15/m0/m18/U3  ( .A(\myram/m15/dout[18] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[18]), .Y(n2155) );
  AOI22X1 \myram/m15/m0/m17/U3  ( .A(\myram/m15/dout[17] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[17]), .Y(n2154) );
  AOI22X1 \myram/m15/m0/m16/U3  ( .A(\myram/m15/dout[16] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[16]), .Y(n2153) );
  AOI22X1 \myram/m15/m0/m15/U3  ( .A(\myram/m15/dout[15] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[15]), .Y(n2152) );
  AOI22X1 \myram/m15/m0/m14/U3  ( .A(\myram/m15/dout[14] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[14]), .Y(n2151) );
  AOI22X1 \myram/m15/m0/m13/U3  ( .A(\myram/m15/dout[13] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[13]), .Y(n2150) );
  AOI22X1 \myram/m15/m0/m12/U3  ( .A(\myram/m15/dout[12] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[12]), .Y(n2149) );
  AOI22X1 \myram/m15/m0/m11/U3  ( .A(\myram/m15/dout[11] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[11]), .Y(n2148) );
  AOI22X1 \myram/m15/m0/m10/U3  ( .A(\myram/m15/dout[10] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[10]), .Y(n2147) );
  AOI22X1 \myram/m15/m0/m9/U3  ( .A(\myram/m15/dout[9] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[9]), .Y(n2146) );
  AOI22X1 \myram/m15/m0/m8/U3  ( .A(\myram/m15/dout[8] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[8]), .Y(n2145) );
  AOI22X1 \myram/m15/m0/m7/U3  ( .A(\myram/m15/dout[7] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[7]), .Y(n2144) );
  AOI22X1 \myram/m15/m0/m6/U3  ( .A(\myram/m15/dout[6] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[6]), .Y(n2143) );
  AOI22X1 \myram/m15/m0/m5/U3  ( .A(\myram/m15/dout[5] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[5]), .Y(n2142) );
  AOI22X1 \myram/m15/m0/m4/U3  ( .A(\myram/m15/dout[4] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[4]), .Y(n2141) );
  AOI22X1 \myram/m15/m0/m3/U3  ( .A(\myram/m15/dout[3] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[3]), .Y(n2140) );
  AOI22X1 \myram/m15/m0/m2/U3  ( .A(\myram/m15/dout[2] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[2]), .Y(n2139) );
  AOI22X1 \myram/m15/m0/m1/U3  ( .A(\myram/m15/dout[1] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[1]), .Y(n2138) );
  AOI22X1 \myram/m15/m0/m0/U3  ( .A(\myram/m15/dout[0] ), .B(n292), .C(
        \myram/sel_s[15] ), .D(mem_s[0]), .Y(n2137) );
  AOI22X1 \myram/m14/m0/m31/U3  ( .A(\myram/m14/dout[31] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(n132), .Y(n2136) );
  AOI22X1 \myram/m14/m0/m30/U3  ( .A(\myram/m14/dout[30] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[30]), .Y(n2135) );
  AOI22X1 \myram/m14/m0/m29/U3  ( .A(\myram/m14/dout[29] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[29]), .Y(n2134) );
  AOI22X1 \myram/m14/m0/m28/U3  ( .A(\myram/m14/dout[28] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[28]), .Y(n2133) );
  AOI22X1 \myram/m14/m0/m27/U3  ( .A(\myram/m14/dout[27] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[27]), .Y(n2132) );
  AOI22X1 \myram/m14/m0/m26/U3  ( .A(\myram/m14/dout[26] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[26]), .Y(n2131) );
  AOI22X1 \myram/m14/m0/m25/U3  ( .A(\myram/m14/dout[25] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[25]), .Y(n2130) );
  AOI22X1 \myram/m14/m0/m24/U3  ( .A(\myram/m14/dout[24] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[24]), .Y(n2129) );
  AOI22X1 \myram/m14/m0/m23/U3  ( .A(\myram/m14/dout[23] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[23]), .Y(n2128) );
  AOI22X1 \myram/m14/m0/m22/U3  ( .A(\myram/m14/dout[22] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[22]), .Y(n2127) );
  AOI22X1 \myram/m14/m0/m21/U3  ( .A(\myram/m14/dout[21] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[21]), .Y(n2126) );
  AOI22X1 \myram/m14/m0/m20/U3  ( .A(\myram/m14/dout[20] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[20]), .Y(n2125) );
  AOI22X1 \myram/m14/m0/m19/U3  ( .A(\myram/m14/dout[19] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[19]), .Y(n2124) );
  AOI22X1 \myram/m14/m0/m18/U3  ( .A(\myram/m14/dout[18] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[18]), .Y(n2123) );
  AOI22X1 \myram/m14/m0/m17/U3  ( .A(\myram/m14/dout[17] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[17]), .Y(n2122) );
  AOI22X1 \myram/m14/m0/m16/U3  ( .A(\myram/m14/dout[16] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[16]), .Y(n2121) );
  AOI22X1 \myram/m14/m0/m15/U3  ( .A(\myram/m14/dout[15] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[15]), .Y(n2120) );
  AOI22X1 \myram/m14/m0/m14/U3  ( .A(\myram/m14/dout[14] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[14]), .Y(n2119) );
  AOI22X1 \myram/m14/m0/m13/U3  ( .A(\myram/m14/dout[13] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[13]), .Y(n2118) );
  AOI22X1 \myram/m14/m0/m12/U3  ( .A(\myram/m14/dout[12] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[12]), .Y(n2117) );
  AOI22X1 \myram/m14/m0/m11/U3  ( .A(\myram/m14/dout[11] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[11]), .Y(n2116) );
  AOI22X1 \myram/m14/m0/m10/U3  ( .A(\myram/m14/dout[10] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[10]), .Y(n2115) );
  AOI22X1 \myram/m14/m0/m9/U3  ( .A(\myram/m14/dout[9] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[9]), .Y(n2114) );
  AOI22X1 \myram/m14/m0/m8/U3  ( .A(\myram/m14/dout[8] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[8]), .Y(n2113) );
  AOI22X1 \myram/m14/m0/m7/U3  ( .A(\myram/m14/dout[7] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[7]), .Y(n2112) );
  AOI22X1 \myram/m14/m0/m6/U3  ( .A(\myram/m14/dout[6] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[6]), .Y(n2111) );
  AOI22X1 \myram/m14/m0/m5/U3  ( .A(\myram/m14/dout[5] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[5]), .Y(n2110) );
  AOI22X1 \myram/m14/m0/m4/U3  ( .A(\myram/m14/dout[4] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[4]), .Y(n2109) );
  AOI22X1 \myram/m14/m0/m3/U3  ( .A(\myram/m14/dout[3] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[3]), .Y(n2108) );
  AOI22X1 \myram/m14/m0/m2/U3  ( .A(\myram/m14/dout[2] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[2]), .Y(n2107) );
  AOI22X1 \myram/m14/m0/m1/U3  ( .A(\myram/m14/dout[1] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[1]), .Y(n2106) );
  AOI22X1 \myram/m14/m0/m0/U3  ( .A(\myram/m14/dout[0] ), .B(n293), .C(
        \myram/sel_s[14] ), .D(mem_s[0]), .Y(n2105) );
  AOI22X1 \myram/m13/m0/m31/U3  ( .A(\myram/m13/dout[31] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(n132), .Y(n2104) );
  AOI22X1 \myram/m13/m0/m30/U3  ( .A(\myram/m13/dout[30] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[30]), .Y(n2103) );
  AOI22X1 \myram/m13/m0/m29/U3  ( .A(\myram/m13/dout[29] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[29]), .Y(n2102) );
  AOI22X1 \myram/m13/m0/m28/U3  ( .A(\myram/m13/dout[28] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[28]), .Y(n2101) );
  AOI22X1 \myram/m13/m0/m27/U3  ( .A(\myram/m13/dout[27] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[27]), .Y(n2100) );
  AOI22X1 \myram/m13/m0/m26/U3  ( .A(\myram/m13/dout[26] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[26]), .Y(n2099) );
  AOI22X1 \myram/m13/m0/m25/U3  ( .A(\myram/m13/dout[25] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[25]), .Y(n2098) );
  AOI22X1 \myram/m13/m0/m24/U3  ( .A(\myram/m13/dout[24] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[24]), .Y(n2097) );
  AOI22X1 \myram/m13/m0/m23/U3  ( .A(\myram/m13/dout[23] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[23]), .Y(n2096) );
  AOI22X1 \myram/m13/m0/m22/U3  ( .A(\myram/m13/dout[22] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[22]), .Y(n2095) );
  AOI22X1 \myram/m13/m0/m21/U3  ( .A(\myram/m13/dout[21] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[21]), .Y(n2094) );
  AOI22X1 \myram/m13/m0/m20/U3  ( .A(\myram/m13/dout[20] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[20]), .Y(n2093) );
  AOI22X1 \myram/m13/m0/m19/U3  ( .A(\myram/m13/dout[19] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[19]), .Y(n2092) );
  AOI22X1 \myram/m13/m0/m18/U3  ( .A(\myram/m13/dout[18] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[18]), .Y(n2091) );
  AOI22X1 \myram/m13/m0/m17/U3  ( .A(\myram/m13/dout[17] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[17]), .Y(n2090) );
  AOI22X1 \myram/m13/m0/m16/U3  ( .A(\myram/m13/dout[16] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[16]), .Y(n2089) );
  AOI22X1 \myram/m13/m0/m15/U3  ( .A(\myram/m13/dout[15] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[15]), .Y(n2088) );
  AOI22X1 \myram/m13/m0/m14/U3  ( .A(\myram/m13/dout[14] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[14]), .Y(n2087) );
  AOI22X1 \myram/m13/m0/m13/U3  ( .A(\myram/m13/dout[13] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[13]), .Y(n2086) );
  AOI22X1 \myram/m13/m0/m12/U3  ( .A(\myram/m13/dout[12] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[12]), .Y(n2085) );
  AOI22X1 \myram/m13/m0/m11/U3  ( .A(\myram/m13/dout[11] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[11]), .Y(n2084) );
  AOI22X1 \myram/m13/m0/m10/U3  ( .A(\myram/m13/dout[10] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[10]), .Y(n2083) );
  AOI22X1 \myram/m13/m0/m9/U3  ( .A(\myram/m13/dout[9] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[9]), .Y(n2082) );
  AOI22X1 \myram/m13/m0/m8/U3  ( .A(\myram/m13/dout[8] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[8]), .Y(n2081) );
  AOI22X1 \myram/m13/m0/m7/U3  ( .A(\myram/m13/dout[7] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[7]), .Y(n2080) );
  AOI22X1 \myram/m13/m0/m6/U3  ( .A(\myram/m13/dout[6] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[6]), .Y(n2079) );
  AOI22X1 \myram/m13/m0/m5/U3  ( .A(\myram/m13/dout[5] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[5]), .Y(n2078) );
  AOI22X1 \myram/m13/m0/m4/U3  ( .A(\myram/m13/dout[4] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[4]), .Y(n2077) );
  AOI22X1 \myram/m13/m0/m3/U3  ( .A(\myram/m13/dout[3] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[3]), .Y(n2076) );
  AOI22X1 \myram/m13/m0/m2/U3  ( .A(\myram/m13/dout[2] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[2]), .Y(n2075) );
  AOI22X1 \myram/m13/m0/m1/U3  ( .A(\myram/m13/dout[1] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[1]), .Y(n2074) );
  AOI22X1 \myram/m13/m0/m0/U3  ( .A(\myram/m13/dout[0] ), .B(n294), .C(
        \myram/sel_s[13] ), .D(mem_s[0]), .Y(n2073) );
  AOI22X1 \myram/m12/m0/m31/U3  ( .A(\myram/m12/dout[31] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(n132), .Y(n2072) );
  AOI22X1 \myram/m12/m0/m30/U3  ( .A(\myram/m12/dout[30] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[30]), .Y(n2071) );
  AOI22X1 \myram/m12/m0/m29/U3  ( .A(\myram/m12/dout[29] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[29]), .Y(n2070) );
  AOI22X1 \myram/m12/m0/m28/U3  ( .A(\myram/m12/dout[28] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[28]), .Y(n2069) );
  AOI22X1 \myram/m12/m0/m27/U3  ( .A(\myram/m12/dout[27] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[27]), .Y(n2068) );
  AOI22X1 \myram/m12/m0/m26/U3  ( .A(\myram/m12/dout[26] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[26]), .Y(n2067) );
  AOI22X1 \myram/m12/m0/m25/U3  ( .A(\myram/m12/dout[25] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[25]), .Y(n2066) );
  AOI22X1 \myram/m12/m0/m24/U3  ( .A(\myram/m12/dout[24] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[24]), .Y(n2065) );
  AOI22X1 \myram/m12/m0/m23/U3  ( .A(\myram/m12/dout[23] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[23]), .Y(n2064) );
  AOI22X1 \myram/m12/m0/m22/U3  ( .A(\myram/m12/dout[22] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[22]), .Y(n2063) );
  AOI22X1 \myram/m12/m0/m21/U3  ( .A(\myram/m12/dout[21] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[21]), .Y(n2062) );
  AOI22X1 \myram/m12/m0/m20/U3  ( .A(\myram/m12/dout[20] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[20]), .Y(n2061) );
  AOI22X1 \myram/m12/m0/m19/U3  ( .A(\myram/m12/dout[19] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[19]), .Y(n2060) );
  AOI22X1 \myram/m12/m0/m18/U3  ( .A(\myram/m12/dout[18] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[18]), .Y(n2059) );
  AOI22X1 \myram/m12/m0/m17/U3  ( .A(\myram/m12/dout[17] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[17]), .Y(n2058) );
  AOI22X1 \myram/m12/m0/m16/U3  ( .A(\myram/m12/dout[16] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[16]), .Y(n2057) );
  AOI22X1 \myram/m12/m0/m15/U3  ( .A(\myram/m12/dout[15] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[15]), .Y(n2056) );
  AOI22X1 \myram/m12/m0/m14/U3  ( .A(\myram/m12/dout[14] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[14]), .Y(n2055) );
  AOI22X1 \myram/m12/m0/m13/U3  ( .A(\myram/m12/dout[13] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[13]), .Y(n2054) );
  AOI22X1 \myram/m12/m0/m12/U3  ( .A(\myram/m12/dout[12] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[12]), .Y(n2053) );
  AOI22X1 \myram/m12/m0/m11/U3  ( .A(\myram/m12/dout[11] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[11]), .Y(n2052) );
  AOI22X1 \myram/m12/m0/m10/U3  ( .A(\myram/m12/dout[10] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[10]), .Y(n2051) );
  AOI22X1 \myram/m12/m0/m9/U3  ( .A(\myram/m12/dout[9] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[9]), .Y(n2050) );
  AOI22X1 \myram/m12/m0/m8/U3  ( .A(\myram/m12/dout[8] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[8]), .Y(n2049) );
  AOI22X1 \myram/m12/m0/m7/U3  ( .A(\myram/m12/dout[7] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[7]), .Y(n2048) );
  AOI22X1 \myram/m12/m0/m6/U3  ( .A(\myram/m12/dout[6] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[6]), .Y(n2047) );
  AOI22X1 \myram/m12/m0/m5/U3  ( .A(\myram/m12/dout[5] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[5]), .Y(n2046) );
  AOI22X1 \myram/m12/m0/m4/U3  ( .A(\myram/m12/dout[4] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[4]), .Y(n2045) );
  AOI22X1 \myram/m12/m0/m3/U3  ( .A(\myram/m12/dout[3] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[3]), .Y(n2044) );
  AOI22X1 \myram/m12/m0/m2/U3  ( .A(\myram/m12/dout[2] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[2]), .Y(n2043) );
  AOI22X1 \myram/m12/m0/m1/U3  ( .A(\myram/m12/dout[1] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[1]), .Y(n2042) );
  AOI22X1 \myram/m12/m0/m0/U3  ( .A(\myram/m12/dout[0] ), .B(n295), .C(
        \myram/sel_s[12] ), .D(mem_s[0]), .Y(n2041) );
  AOI22X1 \myram/m11/m0/m31/U3  ( .A(\myram/m11/dout[31] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(n132), .Y(n2040) );
  AOI22X1 \myram/m11/m0/m30/U3  ( .A(\myram/m11/dout[30] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[30]), .Y(n2039) );
  AOI22X1 \myram/m11/m0/m29/U3  ( .A(\myram/m11/dout[29] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[29]), .Y(n2038) );
  AOI22X1 \myram/m11/m0/m28/U3  ( .A(\myram/m11/dout[28] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[28]), .Y(n2037) );
  AOI22X1 \myram/m11/m0/m27/U3  ( .A(\myram/m11/dout[27] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[27]), .Y(n2036) );
  AOI22X1 \myram/m11/m0/m26/U3  ( .A(\myram/m11/dout[26] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[26]), .Y(n2035) );
  AOI22X1 \myram/m11/m0/m25/U3  ( .A(\myram/m11/dout[25] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[25]), .Y(n2034) );
  AOI22X1 \myram/m11/m0/m24/U3  ( .A(\myram/m11/dout[24] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[24]), .Y(n2033) );
  AOI22X1 \myram/m11/m0/m23/U3  ( .A(\myram/m11/dout[23] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[23]), .Y(n2032) );
  AOI22X1 \myram/m11/m0/m22/U3  ( .A(\myram/m11/dout[22] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[22]), .Y(n2031) );
  AOI22X1 \myram/m11/m0/m21/U3  ( .A(\myram/m11/dout[21] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[21]), .Y(n2030) );
  AOI22X1 \myram/m11/m0/m20/U3  ( .A(\myram/m11/dout[20] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[20]), .Y(n2029) );
  AOI22X1 \myram/m11/m0/m19/U3  ( .A(\myram/m11/dout[19] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[19]), .Y(n2028) );
  AOI22X1 \myram/m11/m0/m18/U3  ( .A(\myram/m11/dout[18] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[18]), .Y(n2027) );
  AOI22X1 \myram/m11/m0/m17/U3  ( .A(\myram/m11/dout[17] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[17]), .Y(n2026) );
  AOI22X1 \myram/m11/m0/m16/U3  ( .A(\myram/m11/dout[16] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[16]), .Y(n2025) );
  AOI22X1 \myram/m11/m0/m15/U3  ( .A(\myram/m11/dout[15] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[15]), .Y(n2024) );
  AOI22X1 \myram/m11/m0/m14/U3  ( .A(\myram/m11/dout[14] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[14]), .Y(n2023) );
  AOI22X1 \myram/m11/m0/m13/U3  ( .A(\myram/m11/dout[13] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[13]), .Y(n2022) );
  AOI22X1 \myram/m11/m0/m12/U3  ( .A(\myram/m11/dout[12] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[12]), .Y(n2021) );
  AOI22X1 \myram/m11/m0/m11/U3  ( .A(\myram/m11/dout[11] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[11]), .Y(n2020) );
  AOI22X1 \myram/m11/m0/m10/U3  ( .A(\myram/m11/dout[10] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[10]), .Y(n2019) );
  AOI22X1 \myram/m11/m0/m9/U3  ( .A(\myram/m11/dout[9] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[9]), .Y(n2018) );
  AOI22X1 \myram/m11/m0/m8/U3  ( .A(\myram/m11/dout[8] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[8]), .Y(n2017) );
  AOI22X1 \myram/m11/m0/m7/U3  ( .A(\myram/m11/dout[7] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[7]), .Y(n2016) );
  AOI22X1 \myram/m11/m0/m6/U3  ( .A(\myram/m11/dout[6] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[6]), .Y(n2015) );
  AOI22X1 \myram/m11/m0/m5/U3  ( .A(\myram/m11/dout[5] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[5]), .Y(n2014) );
  AOI22X1 \myram/m11/m0/m4/U3  ( .A(\myram/m11/dout[4] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[4]), .Y(n2013) );
  AOI22X1 \myram/m11/m0/m3/U3  ( .A(\myram/m11/dout[3] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[3]), .Y(n2012) );
  AOI22X1 \myram/m11/m0/m2/U3  ( .A(\myram/m11/dout[2] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[2]), .Y(n2011) );
  AOI22X1 \myram/m11/m0/m1/U3  ( .A(\myram/m11/dout[1] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[1]), .Y(n2010) );
  AOI22X1 \myram/m11/m0/m0/U3  ( .A(\myram/m11/dout[0] ), .B(n296), .C(
        \myram/sel_s[11] ), .D(mem_s[0]), .Y(n2009) );
  AOI22X1 \myram/m10/m0/m31/U3  ( .A(\myram/m10/dout[31] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[31]), .Y(n2008) );
  AOI22X1 \myram/m10/m0/m30/U3  ( .A(\myram/m10/dout[30] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[30]), .Y(n2007) );
  AOI22X1 \myram/m10/m0/m29/U3  ( .A(\myram/m10/dout[29] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[29]), .Y(n2006) );
  AOI22X1 \myram/m10/m0/m28/U3  ( .A(\myram/m10/dout[28] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[28]), .Y(n2005) );
  AOI22X1 \myram/m10/m0/m27/U3  ( .A(\myram/m10/dout[27] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[27]), .Y(n2004) );
  AOI22X1 \myram/m10/m0/m26/U3  ( .A(\myram/m10/dout[26] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[26]), .Y(n2003) );
  AOI22X1 \myram/m10/m0/m25/U3  ( .A(\myram/m10/dout[25] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[25]), .Y(n2002) );
  AOI22X1 \myram/m10/m0/m24/U3  ( .A(\myram/m10/dout[24] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[24]), .Y(n2001) );
  AOI22X1 \myram/m10/m0/m23/U3  ( .A(\myram/m10/dout[23] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[23]), .Y(n2000) );
  AOI22X1 \myram/m10/m0/m22/U3  ( .A(\myram/m10/dout[22] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[22]), .Y(n1999) );
  AOI22X1 \myram/m10/m0/m21/U3  ( .A(\myram/m10/dout[21] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[21]), .Y(n1998) );
  AOI22X1 \myram/m10/m0/m20/U3  ( .A(\myram/m10/dout[20] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[20]), .Y(n1997) );
  AOI22X1 \myram/m10/m0/m19/U3  ( .A(\myram/m10/dout[19] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[19]), .Y(n1996) );
  AOI22X1 \myram/m10/m0/m18/U3  ( .A(\myram/m10/dout[18] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[18]), .Y(n1995) );
  AOI22X1 \myram/m10/m0/m17/U3  ( .A(\myram/m10/dout[17] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[17]), .Y(n1994) );
  AOI22X1 \myram/m10/m0/m16/U3  ( .A(\myram/m10/dout[16] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[16]), .Y(n1993) );
  AOI22X1 \myram/m10/m0/m15/U3  ( .A(\myram/m10/dout[15] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[15]), .Y(n1992) );
  AOI22X1 \myram/m10/m0/m14/U3  ( .A(\myram/m10/dout[14] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[14]), .Y(n1991) );
  AOI22X1 \myram/m10/m0/m13/U3  ( .A(\myram/m10/dout[13] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[13]), .Y(n1990) );
  AOI22X1 \myram/m10/m0/m12/U3  ( .A(\myram/m10/dout[12] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[12]), .Y(n1989) );
  AOI22X1 \myram/m10/m0/m11/U3  ( .A(\myram/m10/dout[11] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[11]), .Y(n1988) );
  AOI22X1 \myram/m10/m0/m10/U3  ( .A(\myram/m10/dout[10] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[10]), .Y(n1987) );
  AOI22X1 \myram/m10/m0/m9/U3  ( .A(\myram/m10/dout[9] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[9]), .Y(n1986) );
  AOI22X1 \myram/m10/m0/m8/U3  ( .A(\myram/m10/dout[8] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[8]), .Y(n1985) );
  AOI22X1 \myram/m10/m0/m7/U3  ( .A(\myram/m10/dout[7] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[7]), .Y(n1984) );
  AOI22X1 \myram/m10/m0/m6/U3  ( .A(\myram/m10/dout[6] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[6]), .Y(n1983) );
  AOI22X1 \myram/m10/m0/m5/U3  ( .A(\myram/m10/dout[5] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[5]), .Y(n1982) );
  AOI22X1 \myram/m10/m0/m4/U3  ( .A(\myram/m10/dout[4] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[4]), .Y(n1981) );
  AOI22X1 \myram/m10/m0/m3/U3  ( .A(\myram/m10/dout[3] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[3]), .Y(n1980) );
  AOI22X1 \myram/m10/m0/m2/U3  ( .A(\myram/m10/dout[2] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[2]), .Y(n1979) );
  AOI22X1 \myram/m10/m0/m1/U3  ( .A(\myram/m10/dout[1] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[1]), .Y(n1978) );
  AOI22X1 \myram/m10/m0/m0/U3  ( .A(\myram/m10/dout[0] ), .B(n297), .C(
        \myram/sel_s[10] ), .D(mem_s[0]), .Y(n1977) );
  AOI22X1 \myram/m9/m0/m31/U3  ( .A(\myram/m9/dout[31] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(n128), .Y(n1976) );
  AOI22X1 \myram/m9/m0/m30/U3  ( .A(\myram/m9/dout[30] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[30]), .Y(n1975) );
  AOI22X1 \myram/m9/m0/m29/U3  ( .A(\myram/m9/dout[29] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[29]), .Y(n1974) );
  AOI22X1 \myram/m9/m0/m28/U3  ( .A(\myram/m9/dout[28] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[28]), .Y(n1973) );
  AOI22X1 \myram/m9/m0/m27/U3  ( .A(\myram/m9/dout[27] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[27]), .Y(n1972) );
  AOI22X1 \myram/m9/m0/m26/U3  ( .A(\myram/m9/dout[26] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[26]), .Y(n1971) );
  AOI22X1 \myram/m9/m0/m25/U3  ( .A(\myram/m9/dout[25] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[25]), .Y(n1970) );
  AOI22X1 \myram/m9/m0/m24/U3  ( .A(\myram/m9/dout[24] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[24]), .Y(n1969) );
  AOI22X1 \myram/m9/m0/m23/U3  ( .A(\myram/m9/dout[23] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[23]), .Y(n1968) );
  AOI22X1 \myram/m9/m0/m22/U3  ( .A(\myram/m9/dout[22] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[22]), .Y(n1967) );
  AOI22X1 \myram/m9/m0/m21/U3  ( .A(\myram/m9/dout[21] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[21]), .Y(n1966) );
  AOI22X1 \myram/m9/m0/m20/U3  ( .A(\myram/m9/dout[20] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[20]), .Y(n1965) );
  AOI22X1 \myram/m9/m0/m19/U3  ( .A(\myram/m9/dout[19] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[19]), .Y(n1964) );
  AOI22X1 \myram/m9/m0/m18/U3  ( .A(\myram/m9/dout[18] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[18]), .Y(n1963) );
  AOI22X1 \myram/m9/m0/m17/U3  ( .A(\myram/m9/dout[17] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[17]), .Y(n1962) );
  AOI22X1 \myram/m9/m0/m16/U3  ( .A(\myram/m9/dout[16] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[16]), .Y(n1961) );
  AOI22X1 \myram/m9/m0/m15/U3  ( .A(\myram/m9/dout[15] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[15]), .Y(n1960) );
  AOI22X1 \myram/m9/m0/m14/U3  ( .A(\myram/m9/dout[14] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[14]), .Y(n1959) );
  AOI22X1 \myram/m9/m0/m13/U3  ( .A(\myram/m9/dout[13] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[13]), .Y(n1958) );
  AOI22X1 \myram/m9/m0/m12/U3  ( .A(\myram/m9/dout[12] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[12]), .Y(n1957) );
  AOI22X1 \myram/m9/m0/m11/U3  ( .A(\myram/m9/dout[11] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[11]), .Y(n1956) );
  AOI22X1 \myram/m9/m0/m10/U3  ( .A(\myram/m9/dout[10] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[10]), .Y(n1955) );
  AOI22X1 \myram/m9/m0/m9/U3  ( .A(\myram/m9/dout[9] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[9]), .Y(n1954) );
  AOI22X1 \myram/m9/m0/m8/U3  ( .A(\myram/m9/dout[8] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[8]), .Y(n1953) );
  AOI22X1 \myram/m9/m0/m7/U3  ( .A(\myram/m9/dout[7] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[7]), .Y(n1952) );
  AOI22X1 \myram/m9/m0/m6/U3  ( .A(\myram/m9/dout[6] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[6]), .Y(n1951) );
  AOI22X1 \myram/m9/m0/m5/U3  ( .A(\myram/m9/dout[5] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[5]), .Y(n1950) );
  AOI22X1 \myram/m9/m0/m4/U3  ( .A(\myram/m9/dout[4] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[4]), .Y(n1949) );
  AOI22X1 \myram/m9/m0/m3/U3  ( .A(\myram/m9/dout[3] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[3]), .Y(n1948) );
  AOI22X1 \myram/m9/m0/m2/U3  ( .A(\myram/m9/dout[2] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[2]), .Y(n1947) );
  AOI22X1 \myram/m9/m0/m1/U3  ( .A(\myram/m9/dout[1] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[1]), .Y(n1946) );
  AOI22X1 \myram/m9/m0/m0/U3  ( .A(\myram/m9/dout[0] ), .B(n298), .C(
        \myram/sel_s[9] ), .D(mem_s[0]), .Y(n1945) );
  AOI22X1 \myram/m8/m0/m31/U3  ( .A(\myram/m8/dout[31] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[31]), .Y(n1944) );
  AOI22X1 \myram/m8/m0/m30/U3  ( .A(\myram/m8/dout[30] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[30]), .Y(n1943) );
  AOI22X1 \myram/m8/m0/m29/U3  ( .A(\myram/m8/dout[29] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[29]), .Y(n1942) );
  AOI22X1 \myram/m8/m0/m28/U3  ( .A(\myram/m8/dout[28] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[28]), .Y(n1941) );
  AOI22X1 \myram/m8/m0/m27/U3  ( .A(\myram/m8/dout[27] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[27]), .Y(n1940) );
  AOI22X1 \myram/m8/m0/m26/U3  ( .A(\myram/m8/dout[26] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[26]), .Y(n1939) );
  AOI22X1 \myram/m8/m0/m25/U3  ( .A(\myram/m8/dout[25] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[25]), .Y(n1938) );
  AOI22X1 \myram/m8/m0/m24/U3  ( .A(\myram/m8/dout[24] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[24]), .Y(n1937) );
  AOI22X1 \myram/m8/m0/m23/U3  ( .A(\myram/m8/dout[23] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[23]), .Y(n1936) );
  AOI22X1 \myram/m8/m0/m22/U3  ( .A(\myram/m8/dout[22] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[22]), .Y(n1935) );
  AOI22X1 \myram/m8/m0/m21/U3  ( .A(\myram/m8/dout[21] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[21]), .Y(n1934) );
  AOI22X1 \myram/m8/m0/m20/U3  ( .A(\myram/m8/dout[20] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[20]), .Y(n1933) );
  AOI22X1 \myram/m8/m0/m19/U3  ( .A(\myram/m8/dout[19] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[19]), .Y(n1932) );
  AOI22X1 \myram/m8/m0/m18/U3  ( .A(\myram/m8/dout[18] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[18]), .Y(n1931) );
  AOI22X1 \myram/m8/m0/m17/U3  ( .A(\myram/m8/dout[17] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[17]), .Y(n1930) );
  AOI22X1 \myram/m8/m0/m16/U3  ( .A(\myram/m8/dout[16] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[16]), .Y(n1929) );
  AOI22X1 \myram/m8/m0/m15/U3  ( .A(\myram/m8/dout[15] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[15]), .Y(n1928) );
  AOI22X1 \myram/m8/m0/m14/U3  ( .A(\myram/m8/dout[14] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[14]), .Y(n1927) );
  AOI22X1 \myram/m8/m0/m13/U3  ( .A(\myram/m8/dout[13] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[13]), .Y(n1926) );
  AOI22X1 \myram/m8/m0/m12/U3  ( .A(\myram/m8/dout[12] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[12]), .Y(n1925) );
  AOI22X1 \myram/m8/m0/m11/U3  ( .A(\myram/m8/dout[11] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[11]), .Y(n1924) );
  AOI22X1 \myram/m8/m0/m10/U3  ( .A(\myram/m8/dout[10] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[10]), .Y(n1923) );
  AOI22X1 \myram/m8/m0/m9/U3  ( .A(\myram/m8/dout[9] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[9]), .Y(n1922) );
  AOI22X1 \myram/m8/m0/m8/U3  ( .A(\myram/m8/dout[8] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[8]), .Y(n1921) );
  AOI22X1 \myram/m8/m0/m7/U3  ( .A(\myram/m8/dout[7] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[7]), .Y(n1920) );
  AOI22X1 \myram/m8/m0/m6/U3  ( .A(\myram/m8/dout[6] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[6]), .Y(n1919) );
  AOI22X1 \myram/m8/m0/m5/U3  ( .A(\myram/m8/dout[5] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[5]), .Y(n1918) );
  AOI22X1 \myram/m8/m0/m4/U3  ( .A(\myram/m8/dout[4] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[4]), .Y(n1917) );
  AOI22X1 \myram/m8/m0/m3/U3  ( .A(\myram/m8/dout[3] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[3]), .Y(n1916) );
  AOI22X1 \myram/m8/m0/m2/U3  ( .A(\myram/m8/dout[2] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[2]), .Y(n1915) );
  AOI22X1 \myram/m8/m0/m1/U3  ( .A(\myram/m8/dout[1] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[1]), .Y(n1914) );
  AOI22X1 \myram/m8/m0/m0/U3  ( .A(\myram/m8/dout[0] ), .B(n299), .C(
        \myram/sel_s[8] ), .D(mem_s[0]), .Y(n1913) );
  AOI22X1 \myram/m7/m0/m31/U3  ( .A(\myram/m7/dout[31] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(n128), .Y(n1912) );
  AOI22X1 \myram/m7/m0/m30/U3  ( .A(\myram/m7/dout[30] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[30]), .Y(n1911) );
  AOI22X1 \myram/m7/m0/m29/U3  ( .A(\myram/m7/dout[29] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[29]), .Y(n1910) );
  AOI22X1 \myram/m7/m0/m28/U3  ( .A(\myram/m7/dout[28] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[28]), .Y(n1909) );
  AOI22X1 \myram/m7/m0/m27/U3  ( .A(\myram/m7/dout[27] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[27]), .Y(n1908) );
  AOI22X1 \myram/m7/m0/m26/U3  ( .A(\myram/m7/dout[26] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[26]), .Y(n1907) );
  AOI22X1 \myram/m7/m0/m25/U3  ( .A(\myram/m7/dout[25] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[25]), .Y(n1906) );
  AOI22X1 \myram/m7/m0/m24/U3  ( .A(\myram/m7/dout[24] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[24]), .Y(n1905) );
  AOI22X1 \myram/m7/m0/m23/U3  ( .A(\myram/m7/dout[23] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[23]), .Y(n1904) );
  AOI22X1 \myram/m7/m0/m22/U3  ( .A(\myram/m7/dout[22] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[22]), .Y(n1903) );
  AOI22X1 \myram/m7/m0/m21/U3  ( .A(\myram/m7/dout[21] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[21]), .Y(n1902) );
  AOI22X1 \myram/m7/m0/m20/U3  ( .A(\myram/m7/dout[20] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[20]), .Y(n1901) );
  AOI22X1 \myram/m7/m0/m19/U3  ( .A(\myram/m7/dout[19] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[19]), .Y(n1900) );
  AOI22X1 \myram/m7/m0/m18/U3  ( .A(\myram/m7/dout[18] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[18]), .Y(n1899) );
  AOI22X1 \myram/m7/m0/m17/U3  ( .A(\myram/m7/dout[17] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[17]), .Y(n1898) );
  AOI22X1 \myram/m7/m0/m16/U3  ( .A(\myram/m7/dout[16] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[16]), .Y(n1897) );
  AOI22X1 \myram/m7/m0/m15/U3  ( .A(\myram/m7/dout[15] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[15]), .Y(n1896) );
  AOI22X1 \myram/m7/m0/m14/U3  ( .A(\myram/m7/dout[14] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[14]), .Y(n1895) );
  AOI22X1 \myram/m7/m0/m13/U3  ( .A(\myram/m7/dout[13] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[13]), .Y(n1894) );
  AOI22X1 \myram/m7/m0/m12/U3  ( .A(\myram/m7/dout[12] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[12]), .Y(n1893) );
  AOI22X1 \myram/m7/m0/m11/U3  ( .A(\myram/m7/dout[11] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[11]), .Y(n1892) );
  AOI22X1 \myram/m7/m0/m10/U3  ( .A(\myram/m7/dout[10] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[10]), .Y(n1891) );
  AOI22X1 \myram/m7/m0/m9/U3  ( .A(\myram/m7/dout[9] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[9]), .Y(n1890) );
  AOI22X1 \myram/m7/m0/m8/U3  ( .A(\myram/m7/dout[8] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[8]), .Y(n1889) );
  AOI22X1 \myram/m7/m0/m7/U3  ( .A(\myram/m7/dout[7] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[7]), .Y(n1888) );
  AOI22X1 \myram/m7/m0/m6/U3  ( .A(\myram/m7/dout[6] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[6]), .Y(n1887) );
  AOI22X1 \myram/m7/m0/m5/U3  ( .A(\myram/m7/dout[5] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[5]), .Y(n1886) );
  AOI22X1 \myram/m7/m0/m4/U3  ( .A(\myram/m7/dout[4] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[4]), .Y(n1885) );
  AOI22X1 \myram/m7/m0/m3/U3  ( .A(\myram/m7/dout[3] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[3]), .Y(n1884) );
  AOI22X1 \myram/m7/m0/m2/U3  ( .A(\myram/m7/dout[2] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[2]), .Y(n1883) );
  AOI22X1 \myram/m7/m0/m1/U3  ( .A(\myram/m7/dout[1] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[1]), .Y(n1882) );
  AOI22X1 \myram/m7/m0/m0/U3  ( .A(\myram/m7/dout[0] ), .B(n300), .C(
        \myram/sel_s[7] ), .D(mem_s[0]), .Y(n1881) );
  AOI22X1 \myram/m6/m0/m31/U3  ( .A(\myram/m6/dout[31] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[31]), .Y(n1880) );
  AOI22X1 \myram/m6/m0/m30/U3  ( .A(\myram/m6/dout[30] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[30]), .Y(n1879) );
  AOI22X1 \myram/m6/m0/m29/U3  ( .A(\myram/m6/dout[29] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[29]), .Y(n1878) );
  AOI22X1 \myram/m6/m0/m28/U3  ( .A(\myram/m6/dout[28] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[28]), .Y(n1877) );
  AOI22X1 \myram/m6/m0/m27/U3  ( .A(\myram/m6/dout[27] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[27]), .Y(n1876) );
  AOI22X1 \myram/m6/m0/m26/U3  ( .A(\myram/m6/dout[26] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[26]), .Y(n1875) );
  AOI22X1 \myram/m6/m0/m25/U3  ( .A(\myram/m6/dout[25] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[25]), .Y(n1874) );
  AOI22X1 \myram/m6/m0/m24/U3  ( .A(\myram/m6/dout[24] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[24]), .Y(n1873) );
  AOI22X1 \myram/m6/m0/m23/U3  ( .A(\myram/m6/dout[23] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[23]), .Y(n1872) );
  AOI22X1 \myram/m6/m0/m22/U3  ( .A(\myram/m6/dout[22] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[22]), .Y(n1871) );
  AOI22X1 \myram/m6/m0/m21/U3  ( .A(\myram/m6/dout[21] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[21]), .Y(n1870) );
  AOI22X1 \myram/m6/m0/m20/U3  ( .A(\myram/m6/dout[20] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[20]), .Y(n1869) );
  AOI22X1 \myram/m6/m0/m19/U3  ( .A(\myram/m6/dout[19] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[19]), .Y(n1868) );
  AOI22X1 \myram/m6/m0/m18/U3  ( .A(\myram/m6/dout[18] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[18]), .Y(n1867) );
  AOI22X1 \myram/m6/m0/m17/U3  ( .A(\myram/m6/dout[17] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[17]), .Y(n1866) );
  AOI22X1 \myram/m6/m0/m16/U3  ( .A(\myram/m6/dout[16] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[16]), .Y(n1865) );
  AOI22X1 \myram/m6/m0/m15/U3  ( .A(\myram/m6/dout[15] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[15]), .Y(n1864) );
  AOI22X1 \myram/m6/m0/m14/U3  ( .A(\myram/m6/dout[14] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[14]), .Y(n1863) );
  AOI22X1 \myram/m6/m0/m13/U3  ( .A(\myram/m6/dout[13] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[13]), .Y(n1862) );
  AOI22X1 \myram/m6/m0/m12/U3  ( .A(\myram/m6/dout[12] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[12]), .Y(n1861) );
  AOI22X1 \myram/m6/m0/m11/U3  ( .A(\myram/m6/dout[11] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[11]), .Y(n1860) );
  AOI22X1 \myram/m6/m0/m10/U3  ( .A(\myram/m6/dout[10] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[10]), .Y(n1859) );
  AOI22X1 \myram/m6/m0/m9/U3  ( .A(\myram/m6/dout[9] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[9]), .Y(n1858) );
  AOI22X1 \myram/m6/m0/m8/U3  ( .A(\myram/m6/dout[8] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[8]), .Y(n1857) );
  AOI22X1 \myram/m6/m0/m7/U3  ( .A(\myram/m6/dout[7] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[7]), .Y(n1856) );
  AOI22X1 \myram/m6/m0/m6/U3  ( .A(\myram/m6/dout[6] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[6]), .Y(n1855) );
  AOI22X1 \myram/m6/m0/m5/U3  ( .A(\myram/m6/dout[5] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[5]), .Y(n1854) );
  AOI22X1 \myram/m6/m0/m4/U3  ( .A(\myram/m6/dout[4] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[4]), .Y(n1853) );
  AOI22X1 \myram/m6/m0/m3/U3  ( .A(\myram/m6/dout[3] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[3]), .Y(n1852) );
  AOI22X1 \myram/m6/m0/m2/U3  ( .A(\myram/m6/dout[2] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[2]), .Y(n1851) );
  AOI22X1 \myram/m6/m0/m1/U3  ( .A(\myram/m6/dout[1] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[1]), .Y(n1850) );
  AOI22X1 \myram/m6/m0/m0/U3  ( .A(\myram/m6/dout[0] ), .B(n301), .C(
        \myram/sel_s[6] ), .D(mem_s[0]), .Y(n1849) );
  AOI22X1 \myram/m5/m0/m31/U3  ( .A(\myram/m5/dout[31] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(n128), .Y(n1848) );
  AOI22X1 \myram/m5/m0/m30/U3  ( .A(\myram/m5/dout[30] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[30]), .Y(n1847) );
  AOI22X1 \myram/m5/m0/m29/U3  ( .A(\myram/m5/dout[29] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[29]), .Y(n1846) );
  AOI22X1 \myram/m5/m0/m28/U3  ( .A(\myram/m5/dout[28] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[28]), .Y(n1845) );
  AOI22X1 \myram/m5/m0/m27/U3  ( .A(\myram/m5/dout[27] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[27]), .Y(n1844) );
  AOI22X1 \myram/m5/m0/m26/U3  ( .A(\myram/m5/dout[26] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[26]), .Y(n1843) );
  AOI22X1 \myram/m5/m0/m25/U3  ( .A(\myram/m5/dout[25] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[25]), .Y(n1842) );
  AOI22X1 \myram/m5/m0/m24/U3  ( .A(\myram/m5/dout[24] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[24]), .Y(n1841) );
  AOI22X1 \myram/m5/m0/m23/U3  ( .A(\myram/m5/dout[23] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[23]), .Y(n1840) );
  AOI22X1 \myram/m5/m0/m22/U3  ( .A(\myram/m5/dout[22] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[22]), .Y(n1839) );
  AOI22X1 \myram/m5/m0/m21/U3  ( .A(\myram/m5/dout[21] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[21]), .Y(n1838) );
  AOI22X1 \myram/m5/m0/m20/U3  ( .A(\myram/m5/dout[20] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[20]), .Y(n1837) );
  AOI22X1 \myram/m5/m0/m19/U3  ( .A(\myram/m5/dout[19] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[19]), .Y(n1836) );
  AOI22X1 \myram/m5/m0/m18/U3  ( .A(\myram/m5/dout[18] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[18]), .Y(n1835) );
  AOI22X1 \myram/m5/m0/m17/U3  ( .A(\myram/m5/dout[17] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[17]), .Y(n1834) );
  AOI22X1 \myram/m5/m0/m16/U3  ( .A(\myram/m5/dout[16] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[16]), .Y(n1833) );
  AOI22X1 \myram/m5/m0/m15/U3  ( .A(\myram/m5/dout[15] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[15]), .Y(n1832) );
  AOI22X1 \myram/m5/m0/m14/U3  ( .A(\myram/m5/dout[14] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[14]), .Y(n1831) );
  AOI22X1 \myram/m5/m0/m13/U3  ( .A(\myram/m5/dout[13] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[13]), .Y(n1830) );
  AOI22X1 \myram/m5/m0/m12/U3  ( .A(\myram/m5/dout[12] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[12]), .Y(n1829) );
  AOI22X1 \myram/m5/m0/m11/U3  ( .A(\myram/m5/dout[11] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[11]), .Y(n1828) );
  AOI22X1 \myram/m5/m0/m10/U3  ( .A(\myram/m5/dout[10] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[10]), .Y(n1827) );
  AOI22X1 \myram/m5/m0/m9/U3  ( .A(\myram/m5/dout[9] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[9]), .Y(n1826) );
  AOI22X1 \myram/m5/m0/m8/U3  ( .A(\myram/m5/dout[8] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[8]), .Y(n1825) );
  AOI22X1 \myram/m5/m0/m7/U3  ( .A(\myram/m5/dout[7] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[7]), .Y(n1824) );
  AOI22X1 \myram/m5/m0/m6/U3  ( .A(\myram/m5/dout[6] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[6]), .Y(n1823) );
  AOI22X1 \myram/m5/m0/m5/U3  ( .A(\myram/m5/dout[5] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[5]), .Y(n1822) );
  AOI22X1 \myram/m5/m0/m4/U3  ( .A(\myram/m5/dout[4] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[4]), .Y(n1821) );
  AOI22X1 \myram/m5/m0/m3/U3  ( .A(\myram/m5/dout[3] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[3]), .Y(n1820) );
  AOI22X1 \myram/m5/m0/m2/U3  ( .A(\myram/m5/dout[2] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[2]), .Y(n1819) );
  AOI22X1 \myram/m5/m0/m1/U3  ( .A(\myram/m5/dout[1] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[1]), .Y(n1818) );
  AOI22X1 \myram/m5/m0/m0/U3  ( .A(\myram/m5/dout[0] ), .B(n302), .C(
        \myram/sel_s[5] ), .D(mem_s[0]), .Y(n1817) );
  AOI22X1 \myram/m4/m0/m31/U3  ( .A(\myram/m4/dout[31] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[31]), .Y(n1816) );
  AOI22X1 \myram/m4/m0/m30/U3  ( .A(\myram/m4/dout[30] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[30]), .Y(n1815) );
  AOI22X1 \myram/m4/m0/m29/U3  ( .A(\myram/m4/dout[29] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[29]), .Y(n1814) );
  AOI22X1 \myram/m4/m0/m28/U3  ( .A(\myram/m4/dout[28] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[28]), .Y(n1813) );
  AOI22X1 \myram/m4/m0/m27/U3  ( .A(\myram/m4/dout[27] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[27]), .Y(n1812) );
  AOI22X1 \myram/m4/m0/m26/U3  ( .A(\myram/m4/dout[26] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[26]), .Y(n1811) );
  AOI22X1 \myram/m4/m0/m25/U3  ( .A(\myram/m4/dout[25] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[25]), .Y(n1810) );
  AOI22X1 \myram/m4/m0/m24/U3  ( .A(\myram/m4/dout[24] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[24]), .Y(n1809) );
  AOI22X1 \myram/m4/m0/m23/U3  ( .A(\myram/m4/dout[23] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[23]), .Y(n1808) );
  AOI22X1 \myram/m4/m0/m22/U3  ( .A(\myram/m4/dout[22] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[22]), .Y(n1807) );
  AOI22X1 \myram/m4/m0/m21/U3  ( .A(\myram/m4/dout[21] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[21]), .Y(n1806) );
  AOI22X1 \myram/m4/m0/m20/U3  ( .A(\myram/m4/dout[20] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[20]), .Y(n1805) );
  AOI22X1 \myram/m4/m0/m19/U3  ( .A(\myram/m4/dout[19] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[19]), .Y(n1804) );
  AOI22X1 \myram/m4/m0/m18/U3  ( .A(\myram/m4/dout[18] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[18]), .Y(n1803) );
  AOI22X1 \myram/m4/m0/m17/U3  ( .A(\myram/m4/dout[17] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[17]), .Y(n1802) );
  AOI22X1 \myram/m4/m0/m16/U3  ( .A(\myram/m4/dout[16] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[16]), .Y(n1801) );
  AOI22X1 \myram/m4/m0/m15/U3  ( .A(\myram/m4/dout[15] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[15]), .Y(n1800) );
  AOI22X1 \myram/m4/m0/m14/U3  ( .A(\myram/m4/dout[14] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[14]), .Y(n1799) );
  AOI22X1 \myram/m4/m0/m13/U3  ( .A(\myram/m4/dout[13] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[13]), .Y(n1798) );
  AOI22X1 \myram/m4/m0/m12/U3  ( .A(\myram/m4/dout[12] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[12]), .Y(n1797) );
  AOI22X1 \myram/m4/m0/m11/U3  ( .A(\myram/m4/dout[11] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[11]), .Y(n1796) );
  AOI22X1 \myram/m4/m0/m10/U3  ( .A(\myram/m4/dout[10] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[10]), .Y(n1795) );
  AOI22X1 \myram/m4/m0/m9/U3  ( .A(\myram/m4/dout[9] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[9]), .Y(n1794) );
  AOI22X1 \myram/m4/m0/m8/U3  ( .A(\myram/m4/dout[8] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[8]), .Y(n1793) );
  AOI22X1 \myram/m4/m0/m7/U3  ( .A(\myram/m4/dout[7] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[7]), .Y(n1792) );
  AOI22X1 \myram/m4/m0/m6/U3  ( .A(\myram/m4/dout[6] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[6]), .Y(n1791) );
  AOI22X1 \myram/m4/m0/m5/U3  ( .A(\myram/m4/dout[5] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[5]), .Y(n1790) );
  AOI22X1 \myram/m4/m0/m4/U3  ( .A(\myram/m4/dout[4] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[4]), .Y(n1789) );
  AOI22X1 \myram/m4/m0/m3/U3  ( .A(\myram/m4/dout[3] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[3]), .Y(n1788) );
  AOI22X1 \myram/m4/m0/m2/U3  ( .A(\myram/m4/dout[2] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[2]), .Y(n1787) );
  AOI22X1 \myram/m4/m0/m1/U3  ( .A(\myram/m4/dout[1] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[1]), .Y(n1786) );
  AOI22X1 \myram/m4/m0/m0/U3  ( .A(\myram/m4/dout[0] ), .B(n303), .C(
        \myram/sel_s[4] ), .D(mem_s[0]), .Y(n1785) );
  AOI22X1 \myram/m3/m0/m31/U3  ( .A(\myram/m3/dout[31] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(n128), .Y(n1784) );
  AOI22X1 \myram/m3/m0/m30/U3  ( .A(\myram/m3/dout[30] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[30]), .Y(n1783) );
  AOI22X1 \myram/m3/m0/m29/U3  ( .A(\myram/m3/dout[29] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[29]), .Y(n1782) );
  AOI22X1 \myram/m3/m0/m28/U3  ( .A(\myram/m3/dout[28] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[28]), .Y(n1781) );
  AOI22X1 \myram/m3/m0/m27/U3  ( .A(\myram/m3/dout[27] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[27]), .Y(n1780) );
  AOI22X1 \myram/m3/m0/m26/U3  ( .A(\myram/m3/dout[26] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[26]), .Y(n1779) );
  AOI22X1 \myram/m3/m0/m25/U3  ( .A(\myram/m3/dout[25] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[25]), .Y(n1778) );
  AOI22X1 \myram/m3/m0/m24/U3  ( .A(\myram/m3/dout[24] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[24]), .Y(n1777) );
  AOI22X1 \myram/m3/m0/m23/U3  ( .A(\myram/m3/dout[23] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[23]), .Y(n1776) );
  AOI22X1 \myram/m3/m0/m22/U3  ( .A(\myram/m3/dout[22] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[22]), .Y(n1775) );
  AOI22X1 \myram/m3/m0/m21/U3  ( .A(\myram/m3/dout[21] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[21]), .Y(n1774) );
  AOI22X1 \myram/m3/m0/m20/U3  ( .A(\myram/m3/dout[20] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[20]), .Y(n1773) );
  AOI22X1 \myram/m3/m0/m19/U3  ( .A(\myram/m3/dout[19] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[19]), .Y(n1772) );
  AOI22X1 \myram/m3/m0/m18/U3  ( .A(\myram/m3/dout[18] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[18]), .Y(n1771) );
  AOI22X1 \myram/m3/m0/m17/U3  ( .A(\myram/m3/dout[17] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[17]), .Y(n1770) );
  AOI22X1 \myram/m3/m0/m16/U3  ( .A(\myram/m3/dout[16] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[16]), .Y(n1769) );
  AOI22X1 \myram/m3/m0/m15/U3  ( .A(\myram/m3/dout[15] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[15]), .Y(n1768) );
  AOI22X1 \myram/m3/m0/m14/U3  ( .A(\myram/m3/dout[14] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[14]), .Y(n1767) );
  AOI22X1 \myram/m3/m0/m13/U3  ( .A(\myram/m3/dout[13] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[13]), .Y(n1766) );
  AOI22X1 \myram/m3/m0/m12/U3  ( .A(\myram/m3/dout[12] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[12]), .Y(n1765) );
  AOI22X1 \myram/m3/m0/m11/U3  ( .A(\myram/m3/dout[11] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[11]), .Y(n1764) );
  AOI22X1 \myram/m3/m0/m10/U3  ( .A(\myram/m3/dout[10] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[10]), .Y(n1763) );
  AOI22X1 \myram/m3/m0/m9/U3  ( .A(\myram/m3/dout[9] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[9]), .Y(n1762) );
  AOI22X1 \myram/m3/m0/m8/U3  ( .A(\myram/m3/dout[8] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[8]), .Y(n1761) );
  AOI22X1 \myram/m3/m0/m7/U3  ( .A(\myram/m3/dout[7] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[7]), .Y(n1760) );
  AOI22X1 \myram/m3/m0/m6/U3  ( .A(\myram/m3/dout[6] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[6]), .Y(n1759) );
  AOI22X1 \myram/m3/m0/m5/U3  ( .A(\myram/m3/dout[5] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[5]), .Y(n1758) );
  AOI22X1 \myram/m3/m0/m4/U3  ( .A(\myram/m3/dout[4] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[4]), .Y(n1757) );
  AOI22X1 \myram/m3/m0/m3/U3  ( .A(\myram/m3/dout[3] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[3]), .Y(n1756) );
  AOI22X1 \myram/m3/m0/m2/U3  ( .A(\myram/m3/dout[2] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[2]), .Y(n1755) );
  AOI22X1 \myram/m3/m0/m1/U3  ( .A(\myram/m3/dout[1] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[1]), .Y(n1754) );
  AOI22X1 \myram/m3/m0/m0/U3  ( .A(\myram/m3/dout[0] ), .B(n304), .C(
        \myram/sel_s[3] ), .D(mem_s[0]), .Y(n1753) );
  AOI22X1 \myram/m2/m0/m31/U3  ( .A(\myram/m2/dout[31] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[31]), .Y(n1752) );
  AOI22X1 \myram/m2/m0/m30/U3  ( .A(\myram/m2/dout[30] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[30]), .Y(n1751) );
  AOI22X1 \myram/m2/m0/m29/U3  ( .A(\myram/m2/dout[29] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[29]), .Y(n1750) );
  AOI22X1 \myram/m2/m0/m28/U3  ( .A(\myram/m2/dout[28] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[28]), .Y(n1749) );
  AOI22X1 \myram/m2/m0/m27/U3  ( .A(\myram/m2/dout[27] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[27]), .Y(n1748) );
  AOI22X1 \myram/m2/m0/m26/U3  ( .A(\myram/m2/dout[26] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[26]), .Y(n1747) );
  AOI22X1 \myram/m2/m0/m25/U3  ( .A(\myram/m2/dout[25] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[25]), .Y(n1746) );
  AOI22X1 \myram/m2/m0/m24/U3  ( .A(\myram/m2/dout[24] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[24]), .Y(n1745) );
  AOI22X1 \myram/m2/m0/m23/U3  ( .A(\myram/m2/dout[23] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[23]), .Y(n1744) );
  AOI22X1 \myram/m2/m0/m22/U3  ( .A(\myram/m2/dout[22] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[22]), .Y(n1743) );
  AOI22X1 \myram/m2/m0/m21/U3  ( .A(\myram/m2/dout[21] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[21]), .Y(n1742) );
  AOI22X1 \myram/m2/m0/m20/U3  ( .A(\myram/m2/dout[20] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[20]), .Y(n1741) );
  AOI22X1 \myram/m2/m0/m19/U3  ( .A(\myram/m2/dout[19] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[19]), .Y(n1740) );
  AOI22X1 \myram/m2/m0/m18/U3  ( .A(\myram/m2/dout[18] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[18]), .Y(n1739) );
  AOI22X1 \myram/m2/m0/m17/U3  ( .A(\myram/m2/dout[17] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[17]), .Y(n1738) );
  AOI22X1 \myram/m2/m0/m16/U3  ( .A(\myram/m2/dout[16] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[16]), .Y(n1737) );
  AOI22X1 \myram/m2/m0/m15/U3  ( .A(\myram/m2/dout[15] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[15]), .Y(n1736) );
  AOI22X1 \myram/m2/m0/m14/U3  ( .A(\myram/m2/dout[14] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[14]), .Y(n1735) );
  AOI22X1 \myram/m2/m0/m13/U3  ( .A(\myram/m2/dout[13] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[13]), .Y(n1734) );
  AOI22X1 \myram/m2/m0/m12/U3  ( .A(\myram/m2/dout[12] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[12]), .Y(n1733) );
  AOI22X1 \myram/m2/m0/m11/U3  ( .A(\myram/m2/dout[11] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[11]), .Y(n1732) );
  AOI22X1 \myram/m2/m0/m10/U3  ( .A(\myram/m2/dout[10] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[10]), .Y(n1731) );
  AOI22X1 \myram/m2/m0/m9/U3  ( .A(\myram/m2/dout[9] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[9]), .Y(n1730) );
  AOI22X1 \myram/m2/m0/m8/U3  ( .A(\myram/m2/dout[8] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[8]), .Y(n1729) );
  AOI22X1 \myram/m2/m0/m7/U3  ( .A(\myram/m2/dout[7] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[7]), .Y(n1728) );
  AOI22X1 \myram/m2/m0/m6/U3  ( .A(\myram/m2/dout[6] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[6]), .Y(n1727) );
  AOI22X1 \myram/m2/m0/m5/U3  ( .A(\myram/m2/dout[5] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[5]), .Y(n1726) );
  AOI22X1 \myram/m2/m0/m4/U3  ( .A(\myram/m2/dout[4] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[4]), .Y(n1725) );
  AOI22X1 \myram/m2/m0/m3/U3  ( .A(\myram/m2/dout[3] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[3]), .Y(n1724) );
  AOI22X1 \myram/m2/m0/m2/U3  ( .A(\myram/m2/dout[2] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[2]), .Y(n1723) );
  AOI22X1 \myram/m2/m0/m1/U3  ( .A(\myram/m2/dout[1] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[1]), .Y(n1722) );
  AOI22X1 \myram/m2/m0/m0/U3  ( .A(\myram/m2/dout[0] ), .B(n305), .C(
        \myram/sel_s[2] ), .D(mem_s[0]), .Y(n1721) );
  AOI22X1 \myram/m1/m0/m31/U3  ( .A(\myram/m1/dout[31] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(n128), .Y(n1720) );
  AOI22X1 \myram/m1/m0/m30/U3  ( .A(\myram/m1/dout[30] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[30]), .Y(n1719) );
  AOI22X1 \myram/m1/m0/m29/U3  ( .A(\myram/m1/dout[29] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[29]), .Y(n1718) );
  AOI22X1 \myram/m1/m0/m28/U3  ( .A(\myram/m1/dout[28] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[28]), .Y(n1717) );
  AOI22X1 \myram/m1/m0/m27/U3  ( .A(\myram/m1/dout[27] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[27]), .Y(n1716) );
  AOI22X1 \myram/m1/m0/m26/U3  ( .A(\myram/m1/dout[26] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[26]), .Y(n1715) );
  AOI22X1 \myram/m1/m0/m25/U3  ( .A(\myram/m1/dout[25] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[25]), .Y(n1714) );
  AOI22X1 \myram/m1/m0/m24/U3  ( .A(\myram/m1/dout[24] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[24]), .Y(n1713) );
  AOI22X1 \myram/m1/m0/m23/U3  ( .A(\myram/m1/dout[23] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[23]), .Y(n1712) );
  AOI22X1 \myram/m1/m0/m22/U3  ( .A(\myram/m1/dout[22] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[22]), .Y(n1711) );
  AOI22X1 \myram/m1/m0/m21/U3  ( .A(\myram/m1/dout[21] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[21]), .Y(n1710) );
  AOI22X1 \myram/m1/m0/m20/U3  ( .A(\myram/m1/dout[20] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[20]), .Y(n1709) );
  AOI22X1 \myram/m1/m0/m19/U3  ( .A(\myram/m1/dout[19] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[19]), .Y(n1708) );
  AOI22X1 \myram/m1/m0/m18/U3  ( .A(\myram/m1/dout[18] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[18]), .Y(n1707) );
  AOI22X1 \myram/m1/m0/m17/U3  ( .A(\myram/m1/dout[17] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[17]), .Y(n1706) );
  AOI22X1 \myram/m1/m0/m16/U3  ( .A(\myram/m1/dout[16] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[16]), .Y(n1705) );
  AOI22X1 \myram/m1/m0/m15/U3  ( .A(\myram/m1/dout[15] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[15]), .Y(n1704) );
  AOI22X1 \myram/m1/m0/m14/U3  ( .A(\myram/m1/dout[14] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[14]), .Y(n1703) );
  AOI22X1 \myram/m1/m0/m13/U3  ( .A(\myram/m1/dout[13] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[13]), .Y(n1702) );
  AOI22X1 \myram/m1/m0/m12/U3  ( .A(\myram/m1/dout[12] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[12]), .Y(n1701) );
  AOI22X1 \myram/m1/m0/m11/U3  ( .A(\myram/m1/dout[11] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[11]), .Y(n1700) );
  AOI22X1 \myram/m1/m0/m10/U3  ( .A(\myram/m1/dout[10] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[10]), .Y(n1699) );
  AOI22X1 \myram/m1/m0/m9/U3  ( .A(\myram/m1/dout[9] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[9]), .Y(n1698) );
  AOI22X1 \myram/m1/m0/m8/U3  ( .A(\myram/m1/dout[8] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[8]), .Y(n1697) );
  AOI22X1 \myram/m1/m0/m7/U3  ( .A(\myram/m1/dout[7] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[7]), .Y(n1696) );
  AOI22X1 \myram/m1/m0/m6/U3  ( .A(\myram/m1/dout[6] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[6]), .Y(n1695) );
  AOI22X1 \myram/m1/m0/m5/U3  ( .A(\myram/m1/dout[5] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[5]), .Y(n1694) );
  AOI22X1 \myram/m1/m0/m4/U3  ( .A(\myram/m1/dout[4] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[4]), .Y(n1693) );
  AOI22X1 \myram/m1/m0/m3/U3  ( .A(\myram/m1/dout[3] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[3]), .Y(n1692) );
  AOI22X1 \myram/m1/m0/m2/U3  ( .A(\myram/m1/dout[2] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[2]), .Y(n1691) );
  AOI22X1 \myram/m1/m0/m1/U3  ( .A(\myram/m1/dout[1] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[1]), .Y(n1690) );
  AOI22X1 \myram/m1/m0/m0/U3  ( .A(\myram/m1/dout[0] ), .B(n306), .C(
        \myram/sel_s[1] ), .D(mem_s[0]), .Y(n1689) );
  AOI22X1 \myram/m0/m0/m31/U3  ( .A(\myram/m0/dout[31] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[31]), .Y(n1688) );
  AOI22X1 \myram/m0/m0/m30/U3  ( .A(\myram/m0/dout[30] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[30]), .Y(n1687) );
  AOI22X1 \myram/m0/m0/m29/U3  ( .A(\myram/m0/dout[29] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[29]), .Y(n1686) );
  AOI22X1 \myram/m0/m0/m28/U3  ( .A(\myram/m0/dout[28] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[28]), .Y(n1685) );
  AOI22X1 \myram/m0/m0/m27/U3  ( .A(\myram/m0/dout[27] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[27]), .Y(n1684) );
  AOI22X1 \myram/m0/m0/m26/U3  ( .A(\myram/m0/dout[26] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[26]), .Y(n1683) );
  AOI22X1 \myram/m0/m0/m25/U3  ( .A(\myram/m0/dout[25] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[25]), .Y(n1682) );
  AOI22X1 \myram/m0/m0/m24/U3  ( .A(\myram/m0/dout[24] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[24]), .Y(n1681) );
  AOI22X1 \myram/m0/m0/m23/U3  ( .A(\myram/m0/dout[23] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[23]), .Y(n1680) );
  AOI22X1 \myram/m0/m0/m22/U3  ( .A(\myram/m0/dout[22] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[22]), .Y(n1679) );
  AOI22X1 \myram/m0/m0/m21/U3  ( .A(\myram/m0/dout[21] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[21]), .Y(n1678) );
  AOI22X1 \myram/m0/m0/m20/U3  ( .A(\myram/m0/dout[20] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[20]), .Y(n1677) );
  AOI22X1 \myram/m0/m0/m19/U3  ( .A(\myram/m0/dout[19] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[19]), .Y(n1676) );
  AOI22X1 \myram/m0/m0/m18/U3  ( .A(\myram/m0/dout[18] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[18]), .Y(n1675) );
  AOI22X1 \myram/m0/m0/m17/U3  ( .A(\myram/m0/dout[17] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[17]), .Y(n1674) );
  AOI22X1 \myram/m0/m0/m16/U3  ( .A(\myram/m0/dout[16] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[16]), .Y(n1673) );
  AOI22X1 \myram/m0/m0/m15/U3  ( .A(\myram/m0/dout[15] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[15]), .Y(n1672) );
  AOI22X1 \myram/m0/m0/m14/U3  ( .A(\myram/m0/dout[14] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[14]), .Y(n1671) );
  AOI22X1 \myram/m0/m0/m13/U3  ( .A(\myram/m0/dout[13] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[13]), .Y(n1670) );
  AOI22X1 \myram/m0/m0/m12/U3  ( .A(\myram/m0/dout[12] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[12]), .Y(n1669) );
  AOI22X1 \myram/m0/m0/m11/U3  ( .A(\myram/m0/dout[11] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[11]), .Y(n1668) );
  AOI22X1 \myram/m0/m0/m10/U3  ( .A(\myram/m0/dout[10] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[10]), .Y(n1667) );
  AOI22X1 \myram/m0/m0/m9/U3  ( .A(\myram/m0/dout[9] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[9]), .Y(n1666) );
  AOI22X1 \myram/m0/m0/m8/U3  ( .A(\myram/m0/dout[8] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[8]), .Y(n1665) );
  AOI22X1 \myram/m0/m0/m7/U3  ( .A(\myram/m0/dout[7] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[7]), .Y(n1664) );
  AOI22X1 \myram/m0/m0/m6/U3  ( .A(\myram/m0/dout[6] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[6]), .Y(n1663) );
  AOI22X1 \myram/m0/m0/m5/U3  ( .A(\myram/m0/dout[5] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[5]), .Y(n1662) );
  AOI22X1 \myram/m0/m0/m4/U3  ( .A(\myram/m0/dout[4] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[4]), .Y(n1661) );
  AOI22X1 \myram/m0/m0/m3/U3  ( .A(\myram/m0/dout[3] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[3]), .Y(n1660) );
  AOI22X1 \myram/m0/m0/m2/U3  ( .A(\myram/m0/dout[2] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[2]), .Y(n1659) );
  AOI22X1 \myram/m0/m0/m1/U3  ( .A(\myram/m0/dout[1] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[1]), .Y(n1658) );
  AOI22X1 \myram/m0/m0/m0/U3  ( .A(\myram/m0/dout[0] ), .B(n307), .C(
        \myram/sel_s[0] ), .D(mem_s[0]), .Y(n1657) );
  AOI22X1 \myalu/mysrl/mux16/m31/U3  ( .A(\myalu/mysrl/s4[31] ), .B(n1414), 
        .C(b[4]), .D(1'b0), .Y(n1656) );
  AOI22X1 \myalu/mysrl/mux16/m30/U3  ( .A(\myalu/mysrl/s4[30] ), .B(n1624), 
        .C(b[4]), .D(1'b0), .Y(n1655) );
  AOI22X1 \myalu/mysrl/mux16/m29/U3  ( .A(\myalu/mysrl/s4[29] ), .B(n1640), 
        .C(b[4]), .D(1'b0), .Y(n1654) );
  AOI22X1 \myalu/mysrl/mux16/m28/U3  ( .A(\myalu/mysrl/s4[28] ), .B(n1642), 
        .C(b[4]), .D(1'b0), .Y(n1653) );
  AOI22X1 \myalu/mysrl/mux16/m27/U3  ( .A(\myalu/mysrl/s4[27] ), .B(n1650), 
        .C(b[4]), .D(1'b0), .Y(n1652) );
  AOI22X1 \myalu/mysrl/mux16/m26/U3  ( .A(\myalu/mysrl/s4[26] ), .B(n1650), 
        .C(b[4]), .D(1'b0), .Y(n1651) );
  AOI22X1 \myalu/mysrl/mux16/m25/U3  ( .A(\myalu/mysrl/s4[25] ), .B(n1647), 
        .C(b[4]), .D(1'b0), .Y(n1649) );
  AOI22X1 \myalu/mysrl/mux16/m24/U3  ( .A(\myalu/mysrl/s4[24] ), .B(n1647), 
        .C(b[4]), .D(1'b0), .Y(n1648) );
  AOI22X1 \myalu/mysrl/mux16/m23/U3  ( .A(\myalu/mysrl/s4[23] ), .B(n1634), 
        .C(b[4]), .D(1'b0), .Y(n1646) );
  AOI22X1 \myalu/mysrl/mux16/m22/U3  ( .A(\myalu/mysrl/s4[22] ), .B(n1636), 
        .C(b[4]), .D(1'b0), .Y(n1645) );
  AOI22X1 \myalu/mysrl/mux16/m21/U3  ( .A(\myalu/mysrl/s4[21] ), .B(n1638), 
        .C(b[4]), .D(1'b0), .Y(n1644) );
  AOI22X1 \myalu/mysrl/mux16/m20/U3  ( .A(\myalu/mysrl/s4[20] ), .B(n1642), 
        .C(b[4]), .D(1'b0), .Y(n1643) );
  AOI22X1 \myalu/mysrl/mux16/m19/U3  ( .A(\myalu/mysrl/s4[19] ), .B(n1640), 
        .C(b[4]), .D(1'b0), .Y(n1641) );
  AOI22X1 \myalu/mysrl/mux16/m18/U3  ( .A(\myalu/mysrl/s4[18] ), .B(n1638), 
        .C(b[4]), .D(1'b0), .Y(n1639) );
  AOI22X1 \myalu/mysrl/mux16/m17/U3  ( .A(\myalu/mysrl/s4[17] ), .B(n1636), 
        .C(b[4]), .D(1'b0), .Y(n1637) );
  AOI22X1 \myalu/mysrl/mux16/m16/U3  ( .A(\myalu/mysrl/s4[16] ), .B(n1634), 
        .C(b[4]), .D(1'b0), .Y(n1635) );
  AOI22X1 \myalu/mysrl/mux16/m15/U3  ( .A(\myalu/mysrl/s4[15] ), .B(n1622), 
        .C(b[4]), .D(\myalu/mysrl/s4[31] ), .Y(n1633) );
  AOI22X1 \myalu/mysrl/mux16/m14/U3  ( .A(\myalu/mysrl/s4[14] ), .B(n1626), 
        .C(b[4]), .D(\myalu/mysrl/s4[30] ), .Y(n1632) );
  AOI22X1 \myalu/mysrl/mux16/m13/U3  ( .A(\myalu/mysrl/s4[13] ), .B(n1628), 
        .C(b[4]), .D(\myalu/mysrl/s4[29] ), .Y(n1631) );
  AOI22X1 \myalu/mysrl/mux16/m12/U3  ( .A(\myalu/mysrl/s4[12] ), .B(n1370), 
        .C(b[4]), .D(\myalu/mysrl/s4[28] ), .Y(n1630) );
  AOI22X1 \myalu/mysrl/mux16/m11/U3  ( .A(\myalu/mysrl/s4[11] ), .B(n1628), 
        .C(b[4]), .D(\myalu/mysrl/s4[27] ), .Y(n1629) );
  AOI22X1 \myalu/mysrl/mux16/m10/U3  ( .A(\myalu/mysrl/s4[10] ), .B(n1626), 
        .C(b[4]), .D(\myalu/mysrl/s4[26] ), .Y(n1627) );
  AOI22X1 \myalu/mysrl/mux16/m9/U3  ( .A(\myalu/mysrl/s4[9] ), .B(n1624), .C(
        b[4]), .D(\myalu/mysrl/s4[25] ), .Y(n1625) );
  AOI22X1 \myalu/mysrl/mux16/m8/U3  ( .A(\myalu/mysrl/s4[8] ), .B(n1622), .C(
        b[4]), .D(\myalu/mysrl/s4[24] ), .Y(n1623) );
  AOI22X1 \myalu/mysrl/mux16/m7/U3  ( .A(\myalu/mysrl/s4[7] ), .B(n1611), .C(
        b[4]), .D(\myalu/mysrl/s4[23] ), .Y(n1621) );
  AOI22X1 \myalu/mysrl/mux16/m6/U3  ( .A(\myalu/mysrl/s4[6] ), .B(n1613), .C(
        b[4]), .D(\myalu/mysrl/s4[22] ), .Y(n1620) );
  AOI22X1 \myalu/mysrl/mux16/m5/U3  ( .A(\myalu/mysrl/s4[5] ), .B(n1615), .C(
        b[4]), .D(\myalu/mysrl/s4[21] ), .Y(n1619) );
  AOI22X1 \myalu/mysrl/mux16/m4/U3  ( .A(\myalu/mysrl/s4[4] ), .B(n1617), .C(
        b[4]), .D(\myalu/mysrl/s4[20] ), .Y(n1618) );
  AOI22X1 \myalu/mysrl/mux16/m3/U3  ( .A(\myalu/mysrl/s4[3] ), .B(n1615), .C(
        b[4]), .D(\myalu/mysrl/s4[19] ), .Y(n1616) );
  AOI22X1 \myalu/mysrl/mux16/m2/U3  ( .A(\myalu/mysrl/s4[2] ), .B(n1613), .C(
        b[4]), .D(\myalu/mysrl/s4[18] ), .Y(n1614) );
  AOI22X1 \myalu/mysrl/mux16/m1/U3  ( .A(\myalu/mysrl/s4[1] ), .B(n1611), .C(
        b[4]), .D(\myalu/mysrl/s4[17] ), .Y(n1612) );
  AOI22X1 \myalu/mysrl/mux16/m0/U3  ( .A(\myalu/mysrl/s4[0] ), .B(n1609), .C(
        b[4]), .D(\myalu/mysrl/s4[16] ), .Y(n1610) );
  AOI22X1 \myalu/mysrl/mux8/m31/U3  ( .A(\myalu/mysrl/s3[31] ), .B(n1350), .C(
        b[3]), .D(1'b0), .Y(n1608) );
  AOI22X1 \myalu/mysrl/mux8/m30/U3  ( .A(\myalu/mysrl/s3[30] ), .B(n1576), .C(
        b[3]), .D(1'b0), .Y(n1607) );
  AOI22X1 \myalu/mysrl/mux8/m29/U3  ( .A(\myalu/mysrl/s3[29] ), .B(n1604), .C(
        b[3]), .D(1'b0), .Y(n1606) );
  AOI22X1 \myalu/mysrl/mux8/m28/U3  ( .A(\myalu/mysrl/s3[28] ), .B(n1604), .C(
        b[3]), .D(1'b0), .Y(n1605) );
  AOI22X1 \myalu/mysrl/mux8/m27/U3  ( .A(\myalu/mysrl/s3[27] ), .B(n1598), .C(
        b[3]), .D(1'b0), .Y(n1603) );
  AOI22X1 \myalu/mysrl/mux8/m26/U3  ( .A(\myalu/mysrl/s3[26] ), .B(n1600), .C(
        b[3]), .D(1'b0), .Y(n1602) );
  AOI22X1 \myalu/mysrl/mux8/m25/U3  ( .A(\myalu/mysrl/s3[25] ), .B(n1600), .C(
        b[3]), .D(1'b0), .Y(n1601) );
  AOI22X1 \myalu/mysrl/mux8/m24/U3  ( .A(\myalu/mysrl/s3[24] ), .B(n1598), .C(
        b[3]), .D(1'b0), .Y(n1599) );
  AOI22X1 \myalu/mysrl/mux8/m23/U3  ( .A(\myalu/mysrl/s3[23] ), .B(n1589), .C(
        b[3]), .D(\myalu/mysrl/s3[31] ), .Y(n1597) );
  AOI22X1 \myalu/mysrl/mux8/m22/U3  ( .A(\myalu/mysrl/s3[22] ), .B(n1593), .C(
        b[3]), .D(\myalu/mysrl/s3[30] ), .Y(n1596) );
  AOI22X1 \myalu/mysrl/mux8/m21/U3  ( .A(\myalu/mysrl/s3[21] ), .B(n1591), .C(
        b[3]), .D(\myalu/mysrl/s3[29] ), .Y(n1595) );
  AOI22X1 \myalu/mysrl/mux8/m20/U3  ( .A(\myalu/mysrl/s3[20] ), .B(n1593), .C(
        b[3]), .D(\myalu/mysrl/s3[28] ), .Y(n1594) );
  AOI22X1 \myalu/mysrl/mux8/m19/U3  ( .A(\myalu/mysrl/s3[19] ), .B(n1591), .C(
        b[3]), .D(\myalu/mysrl/s3[27] ), .Y(n1592) );
  AOI22X1 \myalu/mysrl/mux8/m18/U3  ( .A(\myalu/mysrl/s3[18] ), .B(n1589), .C(
        b[3]), .D(\myalu/mysrl/s3[26] ), .Y(n1590) );
  AOI22X1 \myalu/mysrl/mux8/m17/U3  ( .A(\myalu/mysrl/s3[17] ), .B(n1574), .C(
        b[3]), .D(\myalu/mysrl/s3[25] ), .Y(n1588) );
  AOI22X1 \myalu/mysrl/mux8/m16/U3  ( .A(\myalu/mysrl/s3[16] ), .B(n1578), .C(
        b[3]), .D(\myalu/mysrl/s3[24] ), .Y(n1587) );
  AOI22X1 \myalu/mysrl/mux8/m15/U3  ( .A(\myalu/mysrl/s3[15] ), .B(n1580), .C(
        b[3]), .D(\myalu/mysrl/s3[23] ), .Y(n1586) );
  AOI22X1 \myalu/mysrl/mux8/m14/U3  ( .A(\myalu/mysrl/s3[14] ), .B(n1582), .C(
        b[3]), .D(\myalu/mysrl/s3[22] ), .Y(n1585) );
  AOI22X1 \myalu/mysrl/mux8/m13/U3  ( .A(\myalu/mysrl/s3[13] ), .B(n1561), .C(
        b[3]), .D(\myalu/mysrl/s3[21] ), .Y(n1584) );
  AOI22X1 \myalu/mysrl/mux8/m12/U3  ( .A(\myalu/mysrl/s3[12] ), .B(n1582), .C(
        b[3]), .D(\myalu/mysrl/s3[20] ), .Y(n1583) );
  AOI22X1 \myalu/mysrl/mux8/m11/U3  ( .A(\myalu/mysrl/s3[11] ), .B(n1580), .C(
        b[3]), .D(\myalu/mysrl/s3[19] ), .Y(n1581) );
  AOI22X1 \myalu/mysrl/mux8/m10/U3  ( .A(\myalu/mysrl/s3[10] ), .B(n1578), .C(
        b[3]), .D(\myalu/mysrl/s3[18] ), .Y(n1579) );
  AOI22X1 \myalu/mysrl/mux8/m9/U3  ( .A(\myalu/mysrl/s3[9] ), .B(n1576), .C(
        b[3]), .D(\myalu/mysrl/s3[17] ), .Y(n1577) );
  AOI22X1 \myalu/mysrl/mux8/m8/U3  ( .A(\myalu/mysrl/s3[8] ), .B(n1574), .C(
        b[3]), .D(\myalu/mysrl/s3[16] ), .Y(n1575) );
  AOI22X1 \myalu/mysrl/mux8/m7/U3  ( .A(\myalu/mysrl/s3[7] ), .B(n1563), .C(
        b[3]), .D(\myalu/mysrl/s3[15] ), .Y(n1573) );
  AOI22X1 \myalu/mysrl/mux8/m6/U3  ( .A(\myalu/mysrl/s3[6] ), .B(n1565), .C(
        b[3]), .D(\myalu/mysrl/s3[14] ), .Y(n1572) );
  AOI22X1 \myalu/mysrl/mux8/m5/U3  ( .A(\myalu/mysrl/s3[5] ), .B(n1567), .C(
        b[3]), .D(\myalu/mysrl/s3[13] ), .Y(n1571) );
  AOI22X1 \myalu/mysrl/mux8/m4/U3  ( .A(\myalu/mysrl/s3[4] ), .B(n1569), .C(
        b[3]), .D(\myalu/mysrl/s3[12] ), .Y(n1570) );
  AOI22X1 \myalu/mysrl/mux8/m3/U3  ( .A(\myalu/mysrl/s3[3] ), .B(n1567), .C(
        b[3]), .D(\myalu/mysrl/s3[11] ), .Y(n1568) );
  AOI22X1 \myalu/mysrl/mux8/m2/U3  ( .A(\myalu/mysrl/s3[2] ), .B(n1565), .C(
        b[3]), .D(\myalu/mysrl/s3[10] ), .Y(n1566) );
  AOI22X1 \myalu/mysrl/mux8/m1/U3  ( .A(\myalu/mysrl/s3[1] ), .B(n1563), .C(
        b[3]), .D(\myalu/mysrl/s3[9] ), .Y(n1564) );
  AOI22X1 \myalu/mysrl/mux8/m0/U3  ( .A(\myalu/mysrl/s3[0] ), .B(n1561), .C(
        b[3]), .D(\myalu/mysrl/s3[8] ), .Y(n1562) );
  AOI22X1 \myalu/mysrl/mux4/m31/U3  ( .A(\myalu/mysrl/s2[31] ), .B(n1286), .C(
        n25), .D(1'b0), .Y(n1560) );
  AOI22X1 \myalu/mysrl/mux4/m30/U3  ( .A(\myalu/mysrl/s2[30] ), .B(n1556), .C(
        n25), .D(1'b0), .Y(n1559) );
  AOI22X1 \myalu/mysrl/mux4/m29/U3  ( .A(\myalu/mysrl/s2[29] ), .B(n1286), .C(
        n25), .D(1'b0), .Y(n1558) );
  AOI22X1 \myalu/mysrl/mux4/m28/U3  ( .A(\myalu/mysrl/s2[28] ), .B(n1556), .C(
        n25), .D(1'b0), .Y(n1557) );
  AOI22X1 \myalu/mysrl/mux4/m27/U3  ( .A(\myalu/mysrl/s2[27] ), .B(n1552), .C(
        n25), .D(\myalu/mysrl/s2[31] ), .Y(n1555) );
  AOI22X1 \myalu/mysrl/mux4/m26/U3  ( .A(\myalu/mysrl/s2[26] ), .B(n1550), .C(
        n25), .D(\myalu/mysrl/s2[30] ), .Y(n1554) );
  AOI22X1 \myalu/mysrl/mux4/m25/U3  ( .A(\myalu/mysrl/s2[25] ), .B(n1552), .C(
        n25), .D(\myalu/mysrl/s2[29] ), .Y(n1553) );
  AOI22X1 \myalu/mysrl/mux4/m24/U3  ( .A(\myalu/mysrl/s2[24] ), .B(n1550), .C(
        n25), .D(\myalu/mysrl/s2[28] ), .Y(n1551) );
  AOI22X1 \myalu/mysrl/mux4/m23/U3  ( .A(\myalu/mysrl/s2[23] ), .B(n1541), .C(
        n25), .D(\myalu/mysrl/s2[27] ), .Y(n1549) );
  AOI22X1 \myalu/mysrl/mux4/m22/U3  ( .A(\myalu/mysrl/s2[22] ), .B(n1545), .C(
        n25), .D(\myalu/mysrl/s2[26] ), .Y(n1548) );
  AOI22X1 \myalu/mysrl/mux4/m21/U3  ( .A(\myalu/mysrl/s2[21] ), .B(n1543), .C(
        n25), .D(\myalu/mysrl/s2[25] ), .Y(n1547) );
  AOI22X1 \myalu/mysrl/mux4/m20/U3  ( .A(\myalu/mysrl/s2[20] ), .B(n1545), .C(
        n25), .D(\myalu/mysrl/s2[24] ), .Y(n1546) );
  AOI22X1 \myalu/mysrl/mux4/m19/U3  ( .A(\myalu/mysrl/s2[19] ), .B(n1543), .C(
        n25), .D(\myalu/mysrl/s2[23] ), .Y(n1544) );
  AOI22X1 \myalu/mysrl/mux4/m18/U3  ( .A(\myalu/mysrl/s2[18] ), .B(n1541), .C(
        n25), .D(\myalu/mysrl/s2[22] ), .Y(n1542) );
  AOI22X1 \myalu/mysrl/mux4/m17/U3  ( .A(\myalu/mysrl/s2[17] ), .B(n1526), .C(
        n25), .D(\myalu/mysrl/s2[21] ), .Y(n1540) );
  AOI22X1 \myalu/mysrl/mux4/m16/U3  ( .A(\myalu/mysrl/s2[16] ), .B(n1528), .C(
        n25), .D(\myalu/mysrl/s2[20] ), .Y(n1539) );
  AOI22X1 \myalu/mysrl/mux4/m15/U3  ( .A(\myalu/mysrl/s2[15] ), .B(n1530), .C(
        n25), .D(\myalu/mysrl/s2[19] ), .Y(n1538) );
  AOI22X1 \myalu/mysrl/mux4/m14/U3  ( .A(\myalu/mysrl/s2[14] ), .B(n1532), .C(
        n25), .D(\myalu/mysrl/s2[18] ), .Y(n1537) );
  AOI22X1 \myalu/mysrl/mux4/m13/U3  ( .A(\myalu/mysrl/s2[13] ), .B(n1534), .C(
        n25), .D(\myalu/mysrl/s2[17] ), .Y(n1536) );
  AOI22X1 \myalu/mysrl/mux4/m12/U3  ( .A(\myalu/mysrl/s2[12] ), .B(n1534), .C(
        n25), .D(\myalu/mysrl/s2[16] ), .Y(n1535) );
  AOI22X1 \myalu/mysrl/mux4/m11/U3  ( .A(\myalu/mysrl/s2[11] ), .B(n1532), .C(
        n25), .D(\myalu/mysrl/s2[15] ), .Y(n1533) );
  AOI22X1 \myalu/mysrl/mux4/m10/U3  ( .A(\myalu/mysrl/s2[10] ), .B(n1530), .C(
        n25), .D(\myalu/mysrl/s2[14] ), .Y(n1531) );
  AOI22X1 \myalu/mysrl/mux4/m9/U3  ( .A(\myalu/mysrl/s2[9] ), .B(n1528), .C(
        n25), .D(\myalu/mysrl/s2[13] ), .Y(n1529) );
  AOI22X1 \myalu/mysrl/mux4/m8/U3  ( .A(\myalu/mysrl/s2[8] ), .B(n1526), .C(
        n25), .D(\myalu/mysrl/s2[12] ), .Y(n1527) );
  AOI22X1 \myalu/mysrl/mux4/m7/U3  ( .A(\myalu/mysrl/s2[7] ), .B(n1515), .C(
        n25), .D(\myalu/mysrl/s2[11] ), .Y(n1525) );
  AOI22X1 \myalu/mysrl/mux4/m6/U3  ( .A(\myalu/mysrl/s2[6] ), .B(n1517), .C(
        n25), .D(\myalu/mysrl/s2[10] ), .Y(n1524) );
  AOI22X1 \myalu/mysrl/mux4/m5/U3  ( .A(\myalu/mysrl/s2[5] ), .B(n1519), .C(
        n25), .D(\myalu/mysrl/s2[9] ), .Y(n1523) );
  AOI22X1 \myalu/mysrl/mux4/m4/U3  ( .A(\myalu/mysrl/s2[4] ), .B(n1521), .C(
        n25), .D(\myalu/mysrl/s2[8] ), .Y(n1522) );
  AOI22X1 \myalu/mysrl/mux4/m3/U3  ( .A(\myalu/mysrl/s2[3] ), .B(n1519), .C(
        n25), .D(\myalu/mysrl/s2[7] ), .Y(n1520) );
  AOI22X1 \myalu/mysrl/mux4/m2/U3  ( .A(\myalu/mysrl/s2[2] ), .B(n1517), .C(
        n25), .D(\myalu/mysrl/s2[6] ), .Y(n1518) );
  AOI22X1 \myalu/mysrl/mux4/m1/U3  ( .A(\myalu/mysrl/s2[1] ), .B(n1515), .C(
        n25), .D(\myalu/mysrl/s2[5] ), .Y(n1516) );
  AOI22X1 \myalu/mysrl/mux4/m0/U3  ( .A(\myalu/mysrl/s2[0] ), .B(n1513), .C(
        n25), .D(\myalu/mysrl/s2[4] ), .Y(n1514) );
  AOI22X1 \myalu/mysrl/mux2/m31/U3  ( .A(\myalu/mysrl/s1[31] ), .B(n1222), .C(
        n62), .D(1'b0), .Y(n1512) );
  AOI22X1 \myalu/mysrl/mux2/m30/U3  ( .A(\myalu/mysrl/s1[30] ), .B(n1509), .C(
        n62), .D(1'b0), .Y(n1511) );
  AOI22X1 \myalu/mysrl/mux2/m29/U3  ( .A(\myalu/mysrl/s1[29] ), .B(n1509), .C(
        n62), .D(\myalu/mysrl/s1[31] ), .Y(n1510) );
  AOI22X1 \myalu/mysrl/mux2/m28/U3  ( .A(\myalu/mysrl/s1[28] ), .B(n1222), .C(
        n62), .D(\myalu/mysrl/s1[30] ), .Y(n1508) );
  AOI22X1 \myalu/mysrl/mux2/m27/U3  ( .A(\myalu/mysrl/s1[27] ), .B(n1504), .C(
        n62), .D(\myalu/mysrl/s1[29] ), .Y(n1507) );
  AOI22X1 \myalu/mysrl/mux2/m26/U3  ( .A(\myalu/mysrl/s1[26] ), .B(n1502), .C(
        n62), .D(\myalu/mysrl/s1[28] ), .Y(n1506) );
  AOI22X1 \myalu/mysrl/mux2/m25/U3  ( .A(\myalu/mysrl/s1[25] ), .B(n1504), .C(
        n62), .D(\myalu/mysrl/s1[27] ), .Y(n1505) );
  AOI22X1 \myalu/mysrl/mux2/m24/U3  ( .A(\myalu/mysrl/s1[24] ), .B(n1502), .C(
        n62), .D(\myalu/mysrl/s1[26] ), .Y(n1503) );
  AOI22X1 \myalu/mysrl/mux2/m23/U3  ( .A(\myalu/mysrl/s1[23] ), .B(n1493), .C(
        n62), .D(\myalu/mysrl/s1[25] ), .Y(n1501) );
  AOI22X1 \myalu/mysrl/mux2/m22/U3  ( .A(\myalu/mysrl/s1[22] ), .B(n1497), .C(
        n62), .D(\myalu/mysrl/s1[24] ), .Y(n1500) );
  AOI22X1 \myalu/mysrl/mux2/m21/U3  ( .A(\myalu/mysrl/s1[21] ), .B(n1495), .C(
        n62), .D(\myalu/mysrl/s1[23] ), .Y(n1499) );
  AOI22X1 \myalu/mysrl/mux2/m20/U3  ( .A(\myalu/mysrl/s1[20] ), .B(n1497), .C(
        n62), .D(\myalu/mysrl/s1[22] ), .Y(n1498) );
  AOI22X1 \myalu/mysrl/mux2/m19/U3  ( .A(\myalu/mysrl/s1[19] ), .B(n1495), .C(
        n62), .D(\myalu/mysrl/s1[21] ), .Y(n1496) );
  AOI22X1 \myalu/mysrl/mux2/m18/U3  ( .A(\myalu/mysrl/s1[18] ), .B(n1493), .C(
        n62), .D(\myalu/mysrl/s1[20] ), .Y(n1494) );
  AOI22X1 \myalu/mysrl/mux2/m17/U3  ( .A(\myalu/mysrl/s1[17] ), .B(n1490), .C(
        n62), .D(\myalu/mysrl/s1[19] ), .Y(n1492) );
  AOI22X1 \myalu/mysrl/mux2/m16/U3  ( .A(\myalu/mysrl/s1[16] ), .B(n1490), .C(
        n62), .D(\myalu/mysrl/s1[18] ), .Y(n1491) );
  AOI22X1 \myalu/mysrl/mux2/m15/U3  ( .A(\myalu/mysrl/s1[15] ), .B(n1479), .C(
        n62), .D(\myalu/mysrl/s1[17] ), .Y(n1489) );
  AOI22X1 \myalu/mysrl/mux2/m14/U3  ( .A(\myalu/mysrl/s1[14] ), .B(n1482), .C(
        n62), .D(\myalu/mysrl/s1[16] ), .Y(n1488) );
  AOI22X1 \myalu/mysrl/mux2/m13/U3  ( .A(\myalu/mysrl/s1[13] ), .B(n1484), .C(
        n62), .D(\myalu/mysrl/s1[15] ), .Y(n1487) );
  AOI22X1 \myalu/mysrl/mux2/m12/U3  ( .A(\myalu/mysrl/s1[12] ), .B(n1467), .C(
        n62), .D(\myalu/mysrl/s1[14] ), .Y(n1486) );
  AOI22X1 \myalu/mysrl/mux2/m11/U3  ( .A(\myalu/mysrl/s1[11] ), .B(n1484), .C(
        n62), .D(\myalu/mysrl/s1[13] ), .Y(n1485) );
  AOI22X1 \myalu/mysrl/mux2/m10/U3  ( .A(\myalu/mysrl/s1[10] ), .B(n1482), .C(
        n62), .D(\myalu/mysrl/s1[12] ), .Y(n1483) );
  AOI22X1 \myalu/mysrl/mux2/m9/U3  ( .A(\myalu/mysrl/s1[9] ), .B(n1465), .C(
        n62), .D(\myalu/mysrl/s1[11] ), .Y(n1481) );
  AOI22X1 \myalu/mysrl/mux2/m8/U3  ( .A(\myalu/mysrl/s1[8] ), .B(n1479), .C(
        n62), .D(\myalu/mysrl/s1[10] ), .Y(n1480) );
  AOI22X1 \myalu/mysrl/mux2/m7/U3  ( .A(\myalu/mysrl/s1[7] ), .B(n1473), .C(
        n62), .D(\myalu/mysrl/s1[9] ), .Y(n1478) );
  AOI22X1 \myalu/mysrl/mux2/m6/U3  ( .A(\myalu/mysrl/s1[6] ), .B(n1475), .C(
        n62), .D(\myalu/mysrl/s1[8] ), .Y(n1477) );
  AOI22X1 \myalu/mysrl/mux2/m5/U3  ( .A(\myalu/mysrl/s1[5] ), .B(n1475), .C(
        n62), .D(\myalu/mysrl/s1[7] ), .Y(n1476) );
  AOI22X1 \myalu/mysrl/mux2/m4/U3  ( .A(\myalu/mysrl/s1[4] ), .B(n1473), .C(
        n62), .D(\myalu/mysrl/s1[6] ), .Y(n1474) );
  AOI22X1 \myalu/mysrl/mux2/m3/U3  ( .A(\myalu/mysrl/s1[3] ), .B(n1471), .C(
        n62), .D(\myalu/mysrl/s1[5] ), .Y(n1472) );
  AOI22X1 \myalu/mysrl/mux2/m2/U3  ( .A(\myalu/mysrl/s1[2] ), .B(n1469), .C(
        n62), .D(\myalu/mysrl/s1[4] ), .Y(n1470) );
  AOI22X1 \myalu/mysrl/mux2/m1/U3  ( .A(\myalu/mysrl/s1[1] ), .B(n1467), .C(
        n62), .D(\myalu/mysrl/s1[3] ), .Y(n1468) );
  AOI22X1 \myalu/mysrl/mux2/m0/U3  ( .A(\myalu/mysrl/s1[0] ), .B(n1465), .C(
        n62), .D(\myalu/mysrl/s1[2] ), .Y(n1466) );
  AOI22X1 \myalu/mysrl/mux1/m31/U3  ( .A(a[31]), .B(n1463), .C(n129), .D(1'b0), 
        .Y(n1464) );
  AOI22X1 \myalu/mysrl/mux1/m30/U3  ( .A(a[30]), .B(n1460), .C(n129), .D(a[31]), .Y(n1462) );
  AOI22X1 \myalu/mysrl/mux1/m29/U3  ( .A(a[29]), .B(n1460), .C(n129), .D(a[30]), .Y(n1461) );
  AOI22X1 \myalu/mysrl/mux1/m28/U3  ( .A(a[28]), .B(n1463), .C(n129), .D(a[29]), .Y(n1459) );
  AOI22X1 \myalu/mysrl/mux1/m27/U3  ( .A(a[27]), .B(n1455), .C(n129), .D(a[28]), .Y(n1458) );
  AOI22X1 \myalu/mysrl/mux1/m26/U3  ( .A(a[26]), .B(n1453), .C(n129), .D(a[27]), .Y(n1457) );
  AOI22X1 \myalu/mysrl/mux1/m25/U3  ( .A(a[25]), .B(n1455), .C(n129), .D(a[26]), .Y(n1456) );
  AOI22X1 \myalu/mysrl/mux1/m24/U3  ( .A(a[24]), .B(n1453), .C(n129), .D(a[25]), .Y(n1454) );
  AOI22X1 \myalu/mysrl/mux1/m23/U3  ( .A(a[23]), .B(n1450), .C(n129), .D(a[24]), .Y(n1452) );
  AOI22X1 \myalu/mysrl/mux1/m22/U3  ( .A(a[22]), .B(n1450), .C(n129), .D(a[23]), .Y(n1451) );
  AOI22X1 \myalu/mysrl/mux1/m21/U3  ( .A(a[21]), .B(n1445), .C(n129), .D(a[22]), .Y(n1449) );
  AOI22X1 \myalu/mysrl/mux1/m20/U3  ( .A(a[20]), .B(n1440), .C(n129), .D(a[21]), .Y(n1448) );
  AOI22X1 \myalu/mysrl/mux1/m19/U3  ( .A(a[19]), .B(n1443), .C(n129), .D(a[20]), .Y(n1447) );
  AOI22X1 \myalu/mysrl/mux1/m18/U3  ( .A(a[18]), .B(n1445), .C(n129), .D(a[19]), .Y(n1446) );
  AOI22X1 \myalu/mysrl/mux1/m17/U3  ( .A(a[17]), .B(n1443), .C(n129), .D(a[18]), .Y(n1444) );
  AOI22X1 \myalu/mysrl/mux1/m16/U3  ( .A(a[16]), .B(n1420), .C(n129), .D(a[17]), .Y(n1442) );
  AOI22X1 \myalu/mysrl/mux1/m15/U3  ( .A(a[15]), .B(n1440), .C(b[0]), .D(a[16]), .Y(n1441) );
  AOI22X1 \myalu/mysrl/mux1/m14/U3  ( .A(a[14]), .B(n1422), .C(n129), .D(a[15]), .Y(n1439) );
  AOI22X1 \myalu/mysrl/mux1/m13/U3  ( .A(a[13]), .B(n1433), .C(b[0]), .D(a[14]), .Y(n1438) );
  AOI22X1 \myalu/mysrl/mux1/m12/U3  ( .A(a[12]), .B(n1435), .C(b[0]), .D(a[13]), .Y(n1437) );
  AOI22X1 \myalu/mysrl/mux1/m11/U3  ( .A(a[11]), .B(n1435), .C(b[0]), .D(a[12]), .Y(n1436) );
  AOI22X1 \myalu/mysrl/mux1/m10/U3  ( .A(a[10]), .B(n1433), .C(b[0]), .D(a[11]), .Y(n1434) );
  AOI22X1 \myalu/mysrl/mux1/m9/U3  ( .A(a[9]), .B(n1418), .C(n129), .D(a[10]), 
        .Y(n1432) );
  AOI22X1 \myalu/mysrl/mux1/m8/U3  ( .A(a[8]), .B(n1157), .C(n129), .D(a[9]), 
        .Y(n1431) );
  AOI22X1 \myalu/mysrl/mux1/m7/U3  ( .A(a[7]), .B(n1424), .C(n129), .D(a[8]), 
        .Y(n1430) );
  AOI22X1 \myalu/mysrl/mux1/m6/U3  ( .A(a[6]), .B(n1428), .C(n129), .D(a[7]), 
        .Y(n1429) );
  AOI22X1 \myalu/mysrl/mux1/m5/U3  ( .A(a[5]), .B(n1426), .C(n129), .D(a[6]), 
        .Y(n1427) );
  AOI22X1 \myalu/mysrl/mux1/m4/U3  ( .A(a[4]), .B(n1424), .C(n129), .D(a[5]), 
        .Y(n1425) );
  AOI22X1 \myalu/mysrl/mux1/m3/U3  ( .A(a[3]), .B(n1422), .C(n129), .D(a[4]), 
        .Y(n1423) );
  AOI22X1 \myalu/mysrl/mux1/m2/U3  ( .A(a[2]), .B(n1420), .C(n129), .D(a[3]), 
        .Y(n1421) );
  AOI22X1 \myalu/mysrl/mux1/m1/U3  ( .A(a[1]), .B(n1418), .C(n129), .D(a[2]), 
        .Y(n1419) );
  AOI22X1 \myalu/mysrl/mux1/m0/U3  ( .A(a[0]), .B(n1416), .C(n129), .D(a[1]), 
        .Y(n1417) );
  AOI22X1 \myalu/mysll/mux16/m31/U3  ( .A(\myalu/mysll/s4[31] ), .B(n1414), 
        .C(b[4]), .D(\myalu/mysll/s4[15] ), .Y(n1415) );
  AOI22X1 \myalu/mysll/mux16/m30/U3  ( .A(\myalu/mysll/s4[30] ), .B(n1412), 
        .C(b[4]), .D(\myalu/mysll/s4[14] ), .Y(n1413) );
  AOI22X1 \myalu/mysll/mux16/m29/U3  ( .A(\myalu/mysll/s4[29] ), .B(n1410), 
        .C(b[4]), .D(\myalu/mysll/s4[13] ), .Y(n1411) );
  AOI22X1 \myalu/mysll/mux16/m28/U3  ( .A(\myalu/mysll/s4[28] ), .B(n1408), 
        .C(b[4]), .D(\myalu/mysll/s4[12] ), .Y(n1409) );
  AOI22X1 \myalu/mysll/mux16/m27/U3  ( .A(\myalu/mysll/s4[27] ), .B(n1406), 
        .C(b[4]), .D(\myalu/mysll/s4[11] ), .Y(n1407) );
  AOI22X1 \myalu/mysll/mux16/m26/U3  ( .A(\myalu/mysll/s4[26] ), .B(n1404), 
        .C(b[4]), .D(\myalu/mysll/s4[10] ), .Y(n1405) );
  AOI22X1 \myalu/mysll/mux16/m25/U3  ( .A(\myalu/mysll/s4[25] ), .B(n1402), 
        .C(b[4]), .D(\myalu/mysll/s4[9] ), .Y(n1403) );
  AOI22X1 \myalu/mysll/mux16/m24/U3  ( .A(\myalu/mysll/s4[24] ), .B(n1400), 
        .C(b[4]), .D(\myalu/mysll/s4[8] ), .Y(n1401) );
  AOI22X1 \myalu/mysll/mux16/m23/U3  ( .A(\myalu/mysll/s4[23] ), .B(n1398), 
        .C(b[4]), .D(\myalu/mysll/s4[7] ), .Y(n1399) );
  AOI22X1 \myalu/mysll/mux16/m22/U3  ( .A(\myalu/mysll/s4[22] ), .B(n1396), 
        .C(b[4]), .D(\myalu/mysll/s4[6] ), .Y(n1397) );
  AOI22X1 \myalu/mysll/mux16/m21/U3  ( .A(\myalu/mysll/s4[21] ), .B(n1394), 
        .C(b[4]), .D(\myalu/mysll/s4[5] ), .Y(n1395) );
  AOI22X1 \myalu/mysll/mux16/m20/U3  ( .A(\myalu/mysll/s4[20] ), .B(n1392), 
        .C(b[4]), .D(\myalu/mysll/s4[4] ), .Y(n1393) );
  AOI22X1 \myalu/mysll/mux16/m19/U3  ( .A(\myalu/mysll/s4[19] ), .B(n1390), 
        .C(b[4]), .D(\myalu/mysll/s4[3] ), .Y(n1391) );
  AOI22X1 \myalu/mysll/mux16/m18/U3  ( .A(\myalu/mysll/s4[18] ), .B(n1388), 
        .C(b[4]), .D(\myalu/mysll/s4[2] ), .Y(n1389) );
  AOI22X1 \myalu/mysll/mux16/m17/U3  ( .A(\myalu/mysll/s4[17] ), .B(n1386), 
        .C(b[4]), .D(\myalu/mysll/s4[1] ), .Y(n1387) );
  AOI22X1 \myalu/mysll/mux16/m16/U3  ( .A(\myalu/mysll/s4[16] ), .B(n1384), 
        .C(b[4]), .D(\myalu/mysll/s4[0] ), .Y(n1385) );
  AOI22X1 \myalu/mysll/mux16/m15/U3  ( .A(\myalu/mysll/s4[15] ), .B(n1382), 
        .C(b[4]), .D(1'b0), .Y(n1383) );
  AOI22X1 \myalu/mysll/mux16/m14/U3  ( .A(\myalu/mysll/s4[14] ), .B(n1380), 
        .C(b[4]), .D(1'b0), .Y(n1381) );
  AOI22X1 \myalu/mysll/mux16/m13/U3  ( .A(\myalu/mysll/s4[13] ), .B(n1378), 
        .C(b[4]), .D(1'b0), .Y(n1379) );
  AOI22X1 \myalu/mysll/mux16/m12/U3  ( .A(\myalu/mysll/s4[12] ), .B(n1376), 
        .C(b[4]), .D(1'b0), .Y(n1377) );
  AOI22X1 \myalu/mysll/mux16/m11/U3  ( .A(\myalu/mysll/s4[11] ), .B(n1374), 
        .C(b[4]), .D(1'b0), .Y(n1375) );
  AOI22X1 \myalu/mysll/mux16/m10/U3  ( .A(\myalu/mysll/s4[10] ), .B(n1372), 
        .C(b[4]), .D(1'b0), .Y(n1373) );
  AOI22X1 \myalu/mysll/mux16/m9/U3  ( .A(\myalu/mysll/s4[9] ), .B(n1370), .C(
        b[4]), .D(1'b0), .Y(n1371) );
  AOI22X1 \myalu/mysll/mux16/m8/U3  ( .A(\myalu/mysll/s4[8] ), .B(n1368), .C(
        b[4]), .D(1'b0), .Y(n1369) );
  AOI22X1 \myalu/mysll/mux16/m7/U3  ( .A(\myalu/mysll/s4[7] ), .B(n1366), .C(
        b[4]), .D(1'b0), .Y(n1367) );
  AOI22X1 \myalu/mysll/mux16/m6/U3  ( .A(\myalu/mysll/s4[6] ), .B(n1364), .C(
        b[4]), .D(1'b0), .Y(n1365) );
  AOI22X1 \myalu/mysll/mux16/m5/U3  ( .A(\myalu/mysll/s4[5] ), .B(n1362), .C(
        b[4]), .D(1'b0), .Y(n1363) );
  AOI22X1 \myalu/mysll/mux16/m4/U3  ( .A(\myalu/mysll/s4[4] ), .B(n1360), .C(
        b[4]), .D(1'b0), .Y(n1361) );
  AOI22X1 \myalu/mysll/mux16/m3/U3  ( .A(\myalu/mysll/s4[3] ), .B(n1358), .C(
        b[4]), .D(1'b0), .Y(n1359) );
  AOI22X1 \myalu/mysll/mux16/m2/U3  ( .A(\myalu/mysll/s4[2] ), .B(n1356), .C(
        b[4]), .D(1'b0), .Y(n1357) );
  AOI22X1 \myalu/mysll/mux16/m1/U3  ( .A(\myalu/mysll/s4[1] ), .B(n1354), .C(
        b[4]), .D(1'b0), .Y(n1355) );
  AOI22X1 \myalu/mysll/mux16/m0/U3  ( .A(\myalu/mysll/s4[0] ), .B(n1352), .C(
        b[4]), .D(1'b0), .Y(n1353) );
  AOI22X1 \myalu/mysll/mux8/m31/U3  ( .A(\myalu/mysll/s3[31] ), .B(n1350), .C(
        b[3]), .D(\myalu/mysll/s3[23] ), .Y(n1351) );
  AOI22X1 \myalu/mysll/mux8/m30/U3  ( .A(\myalu/mysll/s3[30] ), .B(n1348), .C(
        b[3]), .D(\myalu/mysll/s3[22] ), .Y(n1349) );
  AOI22X1 \myalu/mysll/mux8/m29/U3  ( .A(\myalu/mysll/s3[29] ), .B(n1346), .C(
        b[3]), .D(\myalu/mysll/s3[21] ), .Y(n1347) );
  AOI22X1 \myalu/mysll/mux8/m28/U3  ( .A(\myalu/mysll/s3[28] ), .B(n1344), .C(
        b[3]), .D(\myalu/mysll/s3[20] ), .Y(n1345) );
  AOI22X1 \myalu/mysll/mux8/m27/U3  ( .A(\myalu/mysll/s3[27] ), .B(n1342), .C(
        b[3]), .D(\myalu/mysll/s3[19] ), .Y(n1343) );
  AOI22X1 \myalu/mysll/mux8/m26/U3  ( .A(\myalu/mysll/s3[26] ), .B(n1340), .C(
        b[3]), .D(\myalu/mysll/s3[18] ), .Y(n1341) );
  AOI22X1 \myalu/mysll/mux8/m25/U3  ( .A(\myalu/mysll/s3[25] ), .B(n1338), .C(
        b[3]), .D(\myalu/mysll/s3[17] ), .Y(n1339) );
  AOI22X1 \myalu/mysll/mux8/m24/U3  ( .A(\myalu/mysll/s3[24] ), .B(n1336), .C(
        b[3]), .D(\myalu/mysll/s3[16] ), .Y(n1337) );
  AOI22X1 \myalu/mysll/mux8/m23/U3  ( .A(\myalu/mysll/s3[23] ), .B(n1334), .C(
        b[3]), .D(\myalu/mysll/s3[15] ), .Y(n1335) );
  AOI22X1 \myalu/mysll/mux8/m22/U3  ( .A(\myalu/mysll/s3[22] ), .B(n1332), .C(
        b[3]), .D(\myalu/mysll/s3[14] ), .Y(n1333) );
  AOI22X1 \myalu/mysll/mux8/m21/U3  ( .A(\myalu/mysll/s3[21] ), .B(n1330), .C(
        b[3]), .D(\myalu/mysll/s3[13] ), .Y(n1331) );
  AOI22X1 \myalu/mysll/mux8/m20/U3  ( .A(\myalu/mysll/s3[20] ), .B(n1328), .C(
        b[3]), .D(\myalu/mysll/s3[12] ), .Y(n1329) );
  AOI22X1 \myalu/mysll/mux8/m19/U3  ( .A(\myalu/mysll/s3[19] ), .B(n1326), .C(
        b[3]), .D(\myalu/mysll/s3[11] ), .Y(n1327) );
  AOI22X1 \myalu/mysll/mux8/m18/U3  ( .A(\myalu/mysll/s3[18] ), .B(n1324), .C(
        b[3]), .D(\myalu/mysll/s3[10] ), .Y(n1325) );
  AOI22X1 \myalu/mysll/mux8/m17/U3  ( .A(\myalu/mysll/s3[17] ), .B(n1322), .C(
        b[3]), .D(\myalu/mysll/s3[9] ), .Y(n1323) );
  AOI22X1 \myalu/mysll/mux8/m16/U3  ( .A(\myalu/mysll/s3[16] ), .B(n1320), .C(
        b[3]), .D(\myalu/mysll/s3[8] ), .Y(n1321) );
  AOI22X1 \myalu/mysll/mux8/m15/U3  ( .A(\myalu/mysll/s3[15] ), .B(n1318), .C(
        b[3]), .D(\myalu/mysll/s3[7] ), .Y(n1319) );
  AOI22X1 \myalu/mysll/mux8/m14/U3  ( .A(\myalu/mysll/s3[14] ), .B(n1316), .C(
        b[3]), .D(\myalu/mysll/s3[6] ), .Y(n1317) );
  AOI22X1 \myalu/mysll/mux8/m13/U3  ( .A(\myalu/mysll/s3[13] ), .B(n1314), .C(
        b[3]), .D(\myalu/mysll/s3[5] ), .Y(n1315) );
  AOI22X1 \myalu/mysll/mux8/m12/U3  ( .A(\myalu/mysll/s3[12] ), .B(n1312), .C(
        b[3]), .D(\myalu/mysll/s3[4] ), .Y(n1313) );
  AOI22X1 \myalu/mysll/mux8/m11/U3  ( .A(\myalu/mysll/s3[11] ), .B(n1310), .C(
        b[3]), .D(\myalu/mysll/s3[3] ), .Y(n1311) );
  AOI22X1 \myalu/mysll/mux8/m10/U3  ( .A(\myalu/mysll/s3[10] ), .B(n1308), .C(
        b[3]), .D(\myalu/mysll/s3[2] ), .Y(n1309) );
  AOI22X1 \myalu/mysll/mux8/m9/U3  ( .A(\myalu/mysll/s3[9] ), .B(n1306), .C(
        b[3]), .D(\myalu/mysll/s3[1] ), .Y(n1307) );
  AOI22X1 \myalu/mysll/mux8/m8/U3  ( .A(\myalu/mysll/s3[8] ), .B(n1304), .C(
        b[3]), .D(\myalu/mysll/s3[0] ), .Y(n1305) );
  AOI22X1 \myalu/mysll/mux8/m7/U3  ( .A(\myalu/mysll/s3[7] ), .B(n1302), .C(
        b[3]), .D(1'b0), .Y(n1303) );
  AOI22X1 \myalu/mysll/mux8/m6/U3  ( .A(\myalu/mysll/s3[6] ), .B(n1300), .C(
        b[3]), .D(1'b0), .Y(n1301) );
  AOI22X1 \myalu/mysll/mux8/m5/U3  ( .A(\myalu/mysll/s3[5] ), .B(n1298), .C(
        b[3]), .D(1'b0), .Y(n1299) );
  AOI22X1 \myalu/mysll/mux8/m4/U3  ( .A(\myalu/mysll/s3[4] ), .B(n1296), .C(
        b[3]), .D(1'b0), .Y(n1297) );
  AOI22X1 \myalu/mysll/mux8/m3/U3  ( .A(\myalu/mysll/s3[3] ), .B(n1294), .C(
        b[3]), .D(1'b0), .Y(n1295) );
  AOI22X1 \myalu/mysll/mux8/m2/U3  ( .A(\myalu/mysll/s3[2] ), .B(n1292), .C(
        b[3]), .D(1'b0), .Y(n1293) );
  AOI22X1 \myalu/mysll/mux8/m1/U3  ( .A(\myalu/mysll/s3[1] ), .B(n1290), .C(
        b[3]), .D(1'b0), .Y(n1291) );
  AOI22X1 \myalu/mysll/mux8/m0/U3  ( .A(\myalu/mysll/s3[0] ), .B(n1288), .C(
        b[3]), .D(1'b0), .Y(n1289) );
  AOI22X1 \myalu/mysll/mux4/m31/U3  ( .A(\myalu/mysll/s2[31] ), .B(n1286), .C(
        n25), .D(\myalu/mysll/s2[27] ), .Y(n1287) );
  AOI22X1 \myalu/mysll/mux4/m30/U3  ( .A(\myalu/mysll/s2[30] ), .B(n1284), .C(
        n25), .D(\myalu/mysll/s2[26] ), .Y(n1285) );
  AOI22X1 \myalu/mysll/mux4/m29/U3  ( .A(\myalu/mysll/s2[29] ), .B(n1282), .C(
        n25), .D(\myalu/mysll/s2[25] ), .Y(n1283) );
  AOI22X1 \myalu/mysll/mux4/m28/U3  ( .A(\myalu/mysll/s2[28] ), .B(n1280), .C(
        n25), .D(\myalu/mysll/s2[24] ), .Y(n1281) );
  AOI22X1 \myalu/mysll/mux4/m27/U3  ( .A(\myalu/mysll/s2[27] ), .B(n1278), .C(
        n25), .D(\myalu/mysll/s2[23] ), .Y(n1279) );
  AOI22X1 \myalu/mysll/mux4/m26/U3  ( .A(\myalu/mysll/s2[26] ), .B(n1276), .C(
        n25), .D(\myalu/mysll/s2[22] ), .Y(n1277) );
  AOI22X1 \myalu/mysll/mux4/m25/U3  ( .A(\myalu/mysll/s2[25] ), .B(n1274), .C(
        n25), .D(\myalu/mysll/s2[21] ), .Y(n1275) );
  AOI22X1 \myalu/mysll/mux4/m24/U3  ( .A(\myalu/mysll/s2[24] ), .B(n1272), .C(
        n25), .D(\myalu/mysll/s2[20] ), .Y(n1273) );
  AOI22X1 \myalu/mysll/mux4/m23/U3  ( .A(\myalu/mysll/s2[23] ), .B(n1270), .C(
        n25), .D(\myalu/mysll/s2[19] ), .Y(n1271) );
  AOI22X1 \myalu/mysll/mux4/m22/U3  ( .A(\myalu/mysll/s2[22] ), .B(n1268), .C(
        n25), .D(\myalu/mysll/s2[18] ), .Y(n1269) );
  AOI22X1 \myalu/mysll/mux4/m21/U3  ( .A(\myalu/mysll/s2[21] ), .B(n1266), .C(
        n25), .D(\myalu/mysll/s2[17] ), .Y(n1267) );
  AOI22X1 \myalu/mysll/mux4/m20/U3  ( .A(\myalu/mysll/s2[20] ), .B(n1264), .C(
        n25), .D(\myalu/mysll/s2[16] ), .Y(n1265) );
  AOI22X1 \myalu/mysll/mux4/m19/U3  ( .A(\myalu/mysll/s2[19] ), .B(n1262), .C(
        n25), .D(\myalu/mysll/s2[15] ), .Y(n1263) );
  AOI22X1 \myalu/mysll/mux4/m18/U3  ( .A(\myalu/mysll/s2[18] ), .B(n1260), .C(
        n25), .D(\myalu/mysll/s2[14] ), .Y(n1261) );
  AOI22X1 \myalu/mysll/mux4/m17/U3  ( .A(\myalu/mysll/s2[17] ), .B(n1258), .C(
        n25), .D(\myalu/mysll/s2[13] ), .Y(n1259) );
  AOI22X1 \myalu/mysll/mux4/m16/U3  ( .A(\myalu/mysll/s2[16] ), .B(n1256), .C(
        n25), .D(\myalu/mysll/s2[12] ), .Y(n1257) );
  AOI22X1 \myalu/mysll/mux4/m15/U3  ( .A(\myalu/mysll/s2[15] ), .B(n1254), .C(
        n25), .D(\myalu/mysll/s2[11] ), .Y(n1255) );
  AOI22X1 \myalu/mysll/mux4/m14/U3  ( .A(\myalu/mysll/s2[14] ), .B(n1252), .C(
        n25), .D(\myalu/mysll/s2[10] ), .Y(n1253) );
  AOI22X1 \myalu/mysll/mux4/m13/U3  ( .A(\myalu/mysll/s2[13] ), .B(n1250), .C(
        n25), .D(\myalu/mysll/s2[9] ), .Y(n1251) );
  AOI22X1 \myalu/mysll/mux4/m12/U3  ( .A(\myalu/mysll/s2[12] ), .B(n1248), .C(
        n25), .D(\myalu/mysll/s2[8] ), .Y(n1249) );
  AOI22X1 \myalu/mysll/mux4/m11/U3  ( .A(\myalu/mysll/s2[11] ), .B(n1246), .C(
        n25), .D(\myalu/mysll/s2[7] ), .Y(n1247) );
  AOI22X1 \myalu/mysll/mux4/m10/U3  ( .A(\myalu/mysll/s2[10] ), .B(n1244), .C(
        n25), .D(\myalu/mysll/s2[6] ), .Y(n1245) );
  AOI22X1 \myalu/mysll/mux4/m9/U3  ( .A(\myalu/mysll/s2[9] ), .B(n1242), .C(
        n25), .D(\myalu/mysll/s2[5] ), .Y(n1243) );
  AOI22X1 \myalu/mysll/mux4/m8/U3  ( .A(\myalu/mysll/s2[8] ), .B(n1240), .C(
        n25), .D(\myalu/mysll/s2[4] ), .Y(n1241) );
  AOI22X1 \myalu/mysll/mux4/m7/U3  ( .A(\myalu/mysll/s2[7] ), .B(n1238), .C(
        n25), .D(\myalu/mysll/s2[3] ), .Y(n1239) );
  AOI22X1 \myalu/mysll/mux4/m6/U3  ( .A(\myalu/mysll/s2[6] ), .B(n1236), .C(
        n25), .D(\myalu/mysll/s2[2] ), .Y(n1237) );
  AOI22X1 \myalu/mysll/mux4/m5/U3  ( .A(\myalu/mysll/s2[5] ), .B(n1234), .C(
        n25), .D(\myalu/mysll/s2[1] ), .Y(n1235) );
  AOI22X1 \myalu/mysll/mux4/m4/U3  ( .A(\myalu/mysll/s2[4] ), .B(n1232), .C(
        n25), .D(\myalu/mysll/s2[0] ), .Y(n1233) );
  AOI22X1 \myalu/mysll/mux4/m3/U3  ( .A(\myalu/mysll/s2[3] ), .B(n1230), .C(
        n25), .D(1'b0), .Y(n1231) );
  AOI22X1 \myalu/mysll/mux4/m2/U3  ( .A(\myalu/mysll/s2[2] ), .B(n1228), .C(
        n25), .D(1'b0), .Y(n1229) );
  AOI22X1 \myalu/mysll/mux4/m1/U3  ( .A(\myalu/mysll/s2[1] ), .B(n1226), .C(
        n25), .D(1'b0), .Y(n1227) );
  AOI22X1 \myalu/mysll/mux4/m0/U3  ( .A(\myalu/mysll/s2[0] ), .B(n1224), .C(
        n25), .D(1'b0), .Y(n1225) );
  AOI22X1 \myalu/mysll/mux2/m31/U3  ( .A(\myalu/mysll/s1[31] ), .B(n1222), .C(
        n62), .D(\myalu/mysll/s1[29] ), .Y(n1223) );
  AOI22X1 \myalu/mysll/mux2/m30/U3  ( .A(\myalu/mysll/s1[30] ), .B(n1220), .C(
        n62), .D(\myalu/mysll/s1[28] ), .Y(n1221) );
  AOI22X1 \myalu/mysll/mux2/m29/U3  ( .A(\myalu/mysll/s1[29] ), .B(n1218), .C(
        n62), .D(\myalu/mysll/s1[27] ), .Y(n1219) );
  AOI22X1 \myalu/mysll/mux2/m28/U3  ( .A(\myalu/mysll/s1[28] ), .B(n1216), .C(
        n62), .D(\myalu/mysll/s1[26] ), .Y(n1217) );
  AOI22X1 \myalu/mysll/mux2/m27/U3  ( .A(\myalu/mysll/s1[27] ), .B(n1214), .C(
        n62), .D(\myalu/mysll/s1[25] ), .Y(n1215) );
  AOI22X1 \myalu/mysll/mux2/m26/U3  ( .A(\myalu/mysll/s1[26] ), .B(n1212), .C(
        n62), .D(\myalu/mysll/s1[24] ), .Y(n1213) );
  AOI22X1 \myalu/mysll/mux2/m25/U3  ( .A(\myalu/mysll/s1[25] ), .B(n1210), .C(
        n62), .D(\myalu/mysll/s1[23] ), .Y(n1211) );
  AOI22X1 \myalu/mysll/mux2/m24/U3  ( .A(\myalu/mysll/s1[24] ), .B(n1208), .C(
        n62), .D(\myalu/mysll/s1[22] ), .Y(n1209) );
  AOI22X1 \myalu/mysll/mux2/m23/U3  ( .A(\myalu/mysll/s1[23] ), .B(n1206), .C(
        n62), .D(\myalu/mysll/s1[21] ), .Y(n1207) );
  AOI22X1 \myalu/mysll/mux2/m22/U3  ( .A(\myalu/mysll/s1[22] ), .B(n1204), .C(
        n62), .D(\myalu/mysll/s1[20] ), .Y(n1205) );
  AOI22X1 \myalu/mysll/mux2/m21/U3  ( .A(\myalu/mysll/s1[21] ), .B(n1202), .C(
        n62), .D(\myalu/mysll/s1[19] ), .Y(n1203) );
  AOI22X1 \myalu/mysll/mux2/m20/U3  ( .A(\myalu/mysll/s1[20] ), .B(n1200), .C(
        n62), .D(\myalu/mysll/s1[18] ), .Y(n1201) );
  AOI22X1 \myalu/mysll/mux2/m19/U3  ( .A(\myalu/mysll/s1[19] ), .B(n1198), .C(
        n62), .D(\myalu/mysll/s1[17] ), .Y(n1199) );
  AOI22X1 \myalu/mysll/mux2/m18/U3  ( .A(\myalu/mysll/s1[18] ), .B(n1196), .C(
        n62), .D(\myalu/mysll/s1[16] ), .Y(n1197) );
  AOI22X1 \myalu/mysll/mux2/m17/U3  ( .A(\myalu/mysll/s1[17] ), .B(n1194), .C(
        n62), .D(\myalu/mysll/s1[15] ), .Y(n1195) );
  AOI22X1 \myalu/mysll/mux2/m16/U3  ( .A(\myalu/mysll/s1[16] ), .B(n1192), .C(
        n62), .D(\myalu/mysll/s1[14] ), .Y(n1193) );
  AOI22X1 \myalu/mysll/mux2/m15/U3  ( .A(\myalu/mysll/s1[15] ), .B(n1190), .C(
        n62), .D(\myalu/mysll/s1[13] ), .Y(n1191) );
  AOI22X1 \myalu/mysll/mux2/m14/U3  ( .A(\myalu/mysll/s1[14] ), .B(n1188), .C(
        n62), .D(\myalu/mysll/s1[12] ), .Y(n1189) );
  AOI22X1 \myalu/mysll/mux2/m13/U3  ( .A(\myalu/mysll/s1[13] ), .B(n1186), .C(
        n62), .D(\myalu/mysll/s1[11] ), .Y(n1187) );
  AOI22X1 \myalu/mysll/mux2/m12/U3  ( .A(\myalu/mysll/s1[12] ), .B(n1184), .C(
        n62), .D(\myalu/mysll/s1[10] ), .Y(n1185) );
  AOI22X1 \myalu/mysll/mux2/m11/U3  ( .A(\myalu/mysll/s1[11] ), .B(n1182), .C(
        n62), .D(\myalu/mysll/s1[9] ), .Y(n1183) );
  AOI22X1 \myalu/mysll/mux2/m10/U3  ( .A(\myalu/mysll/s1[10] ), .B(n1180), .C(
        n62), .D(\myalu/mysll/s1[8] ), .Y(n1181) );
  AOI22X1 \myalu/mysll/mux2/m9/U3  ( .A(\myalu/mysll/s1[9] ), .B(n1178), .C(
        n62), .D(\myalu/mysll/s1[7] ), .Y(n1179) );
  AOI22X1 \myalu/mysll/mux2/m8/U3  ( .A(\myalu/mysll/s1[8] ), .B(n1176), .C(
        n62), .D(\myalu/mysll/s1[6] ), .Y(n1177) );
  AOI22X1 \myalu/mysll/mux2/m7/U3  ( .A(\myalu/mysll/s1[7] ), .B(n1174), .C(
        n62), .D(\myalu/mysll/s1[5] ), .Y(n1175) );
  AOI22X1 \myalu/mysll/mux2/m6/U3  ( .A(\myalu/mysll/s1[6] ), .B(n1172), .C(
        n62), .D(\myalu/mysll/s1[4] ), .Y(n1173) );
  AOI22X1 \myalu/mysll/mux2/m5/U3  ( .A(\myalu/mysll/s1[5] ), .B(n1170), .C(
        n62), .D(\myalu/mysll/s1[3] ), .Y(n1171) );
  AOI22X1 \myalu/mysll/mux2/m4/U3  ( .A(\myalu/mysll/s1[4] ), .B(n1168), .C(
        n62), .D(\myalu/mysll/s1[2] ), .Y(n1169) );
  AOI22X1 \myalu/mysll/mux2/m3/U3  ( .A(\myalu/mysll/s1[3] ), .B(n1166), .C(
        n62), .D(\myalu/mysll/s1[1] ), .Y(n1167) );
  AOI22X1 \myalu/mysll/mux2/m2/U3  ( .A(\myalu/mysll/s1[2] ), .B(n1164), .C(
        n62), .D(\myalu/mysll/s1[0] ), .Y(n1165) );
  AOI22X1 \myalu/mysll/mux2/m1/U3  ( .A(\myalu/mysll/s1[1] ), .B(n1162), .C(
        n62), .D(1'b0), .Y(n1163) );
  AOI22X1 \myalu/mysll/mux2/m0/U3  ( .A(\myalu/mysll/s1[0] ), .B(n1160), .C(
        n62), .D(1'b0), .Y(n1161) );
  AOI22X1 \myalu/mysll/mux1/m31/U3  ( .A(a[31]), .B(n1463), .C(n129), .D(a[30]), .Y(n1159) );
  AOI22X1 \myalu/mysll/mux1/m30/U3  ( .A(a[30]), .B(n1157), .C(n129), .D(a[29]), .Y(n1158) );
  AOI22X1 \myalu/mysll/mux1/m29/U3  ( .A(a[29]), .B(n1155), .C(n129), .D(a[28]), .Y(n1156) );
  AOI22X1 \myalu/mysll/mux1/m28/U3  ( .A(a[28]), .B(n1153), .C(n129), .D(a[27]), .Y(n1154) );
  AOI22X1 \myalu/mysll/mux1/m27/U3  ( .A(a[27]), .B(n1151), .C(b[0]), .D(a[26]), .Y(n1152) );
  AOI22X1 \myalu/mysll/mux1/m26/U3  ( .A(a[26]), .B(n1149), .C(b[0]), .D(a[25]), .Y(n1150) );
  AOI22X1 \myalu/mysll/mux1/m25/U3  ( .A(a[25]), .B(n1147), .C(b[0]), .D(a[24]), .Y(n1148) );
  AOI22X1 \myalu/mysll/mux1/m24/U3  ( .A(a[24]), .B(n1145), .C(b[0]), .D(a[23]), .Y(n1146) );
  AOI22X1 \myalu/mysll/mux1/m23/U3  ( .A(a[23]), .B(n1143), .C(b[0]), .D(a[22]), .Y(n1144) );
  AOI22X1 \myalu/mysll/mux1/m22/U3  ( .A(a[22]), .B(n1141), .C(b[0]), .D(a[21]), .Y(n1142) );
  AOI22X1 \myalu/mysll/mux1/m21/U3  ( .A(a[21]), .B(n1139), .C(b[0]), .D(a[20]), .Y(n1140) );
  AOI22X1 \myalu/mysll/mux1/m20/U3  ( .A(a[20]), .B(n1137), .C(b[0]), .D(a[19]), .Y(n1138) );
  AOI22X1 \myalu/mysll/mux1/m19/U3  ( .A(a[19]), .B(n1135), .C(b[0]), .D(a[18]), .Y(n1136) );
  AOI22X1 \myalu/mysll/mux1/m18/U3  ( .A(a[18]), .B(n1133), .C(b[0]), .D(a[17]), .Y(n1134) );
  AOI22X1 \myalu/mysll/mux1/m17/U3  ( .A(a[17]), .B(n1131), .C(b[0]), .D(a[16]), .Y(n1132) );
  AOI22X1 \myalu/mysll/mux1/m16/U3  ( .A(a[16]), .B(n1129), .C(b[0]), .D(a[15]), .Y(n1130) );
  AOI22X1 \myalu/mysll/mux1/m15/U3  ( .A(a[15]), .B(n1127), .C(b[0]), .D(a[14]), .Y(n1128) );
  AOI22X1 \myalu/mysll/mux1/m14/U3  ( .A(a[14]), .B(n1125), .C(b[0]), .D(a[13]), .Y(n1126) );
  AOI22X1 \myalu/mysll/mux1/m13/U3  ( .A(a[13]), .B(n1123), .C(b[0]), .D(a[12]), .Y(n1124) );
  AOI22X1 \myalu/mysll/mux1/m12/U3  ( .A(a[12]), .B(n1121), .C(b[0]), .D(a[11]), .Y(n1122) );
  AOI22X1 \myalu/mysll/mux1/m11/U3  ( .A(a[11]), .B(n1119), .C(b[0]), .D(a[10]), .Y(n1120) );
  AOI22X1 \myalu/mysll/mux1/m10/U3  ( .A(a[10]), .B(n1117), .C(b[0]), .D(a[9]), 
        .Y(n1118) );
  AOI22X1 \myalu/mysll/mux1/m9/U3  ( .A(a[9]), .B(n1115), .C(b[0]), .D(a[8]), 
        .Y(n1116) );
  AOI22X1 \myalu/mysll/mux1/m8/U3  ( .A(a[8]), .B(n1113), .C(b[0]), .D(a[7]), 
        .Y(n1114) );
  AOI22X1 \myalu/mysll/mux1/m7/U3  ( .A(a[7]), .B(n1111), .C(n129), .D(a[6]), 
        .Y(n1112) );
  AOI22X1 \myalu/mysll/mux1/m6/U3  ( .A(a[6]), .B(n1109), .C(n129), .D(a[5]), 
        .Y(n1110) );
  AOI22X1 \myalu/mysll/mux1/m5/U3  ( .A(a[5]), .B(n1107), .C(n129), .D(a[4]), 
        .Y(n1108) );
  AOI22X1 \myalu/mysll/mux1/m4/U3  ( .A(a[4]), .B(n1105), .C(n129), .D(a[3]), 
        .Y(n1106) );
  AOI22X1 \myalu/mysll/mux1/m3/U3  ( .A(a[3]), .B(n1103), .C(n129), .D(a[2]), 
        .Y(n1104) );
  AOI22X1 \myalu/mysll/mux1/m2/U3  ( .A(a[2]), .B(n1101), .C(n129), .D(a[1]), 
        .Y(n1102) );
  AOI22X1 \myalu/mysll/mux1/m1/U3  ( .A(a[1]), .B(n1099), .C(n129), .D(a[0]), 
        .Y(n1100) );
  AOI22X1 \myalu/mysll/mux1/m0/U3  ( .A(a[0]), .B(n1097), .C(n129), .D(1'b0), 
        .Y(n1098) );
  AOI22X1 \myalu/muxs/m31/U3  ( .A(\myalu/s0[31] ), .B(n314), .C(alu_op[2]), 
        .D(n185), .Y(n1096) );
  AOI22X1 \myalu/muxs/m30/U3  ( .A(\myalu/s0[30] ), .B(n314), .C(alu_op[2]), 
        .D(n183), .Y(n1095) );
  AOI22X1 \myalu/muxs/m29/U3  ( .A(\myalu/s0[29] ), .B(n314), .C(alu_op[2]), 
        .D(n182), .Y(n1094) );
  AOI22X1 \myalu/muxs/m28/U3  ( .A(\myalu/s0[28] ), .B(n314), .C(alu_op[2]), 
        .D(n181), .Y(n1093) );
  AOI22X1 \myalu/muxs/m27/U3  ( .A(\myalu/s0[27] ), .B(n314), .C(alu_op[2]), 
        .D(n180), .Y(n1092) );
  AOI22X1 \myalu/muxs/m26/U3  ( .A(\myalu/s0[26] ), .B(n314), .C(alu_op[2]), 
        .D(n179), .Y(n1091) );
  AOI22X1 \myalu/muxs/m25/U3  ( .A(\myalu/s0[25] ), .B(n314), .C(alu_op[2]), 
        .D(n178), .Y(n1090) );
  AOI22X1 \myalu/muxs/m24/U3  ( .A(\myalu/s0[24] ), .B(n314), .C(alu_op[2]), 
        .D(n177), .Y(n1089) );
  AOI22X1 \myalu/muxs/m23/U3  ( .A(\myalu/s0[23] ), .B(n314), .C(alu_op[2]), 
        .D(n176), .Y(n1088) );
  AOI22X1 \myalu/muxs/m22/U3  ( .A(\myalu/s0[22] ), .B(n314), .C(alu_op[2]), 
        .D(n175), .Y(n1087) );
  AOI22X1 \myalu/muxs/m21/U3  ( .A(\myalu/s0[21] ), .B(n314), .C(alu_op[2]), 
        .D(n174), .Y(n1086) );
  AOI22X1 \myalu/muxs/m20/U3  ( .A(\myalu/s0[20] ), .B(n314), .C(alu_op[2]), 
        .D(n173), .Y(n1085) );
  AOI22X1 \myalu/muxs/m19/U3  ( .A(\myalu/s0[19] ), .B(n314), .C(alu_op[2]), 
        .D(n172), .Y(n1084) );
  AOI22X1 \myalu/muxs/m18/U3  ( .A(\myalu/s0[18] ), .B(n314), .C(alu_op[2]), 
        .D(n171), .Y(n1083) );
  AOI22X1 \myalu/muxs/m17/U3  ( .A(\myalu/s0[17] ), .B(n314), .C(alu_op[2]), 
        .D(n170), .Y(n1082) );
  AOI22X1 \myalu/muxs/m16/U3  ( .A(\myalu/s0[16] ), .B(n314), .C(alu_op[2]), 
        .D(n154), .Y(n1081) );
  AOI22X1 \myalu/muxs/m15/U3  ( .A(\myalu/s0[15] ), .B(n314), .C(alu_op[2]), 
        .D(n168), .Y(n1080) );
  AOI22X1 \myalu/muxs/m14/U3  ( .A(\myalu/s0[14] ), .B(n314), .C(alu_op[2]), 
        .D(n167), .Y(n1079) );
  AOI22X1 \myalu/muxs/m13/U3  ( .A(\myalu/s0[13] ), .B(n314), .C(alu_op[2]), 
        .D(n166), .Y(n1078) );
  AOI22X1 \myalu/muxs/m12/U3  ( .A(\myalu/s0[12] ), .B(n314), .C(alu_op[2]), 
        .D(n165), .Y(n1077) );
  AOI22X1 \myalu/muxs/m11/U3  ( .A(\myalu/s0[11] ), .B(n314), .C(alu_op[2]), 
        .D(n164), .Y(n1076) );
  AOI22X1 \myalu/muxs/m10/U3  ( .A(\myalu/s0[10] ), .B(n314), .C(alu_op[2]), 
        .D(n163), .Y(n1075) );
  AOI22X1 \myalu/muxs/m9/U3  ( .A(\myalu/s0[9] ), .B(n314), .C(alu_op[2]), .D(
        n153), .Y(n1074) );
  AOI22X1 \myalu/muxs/m8/U3  ( .A(\myalu/s0[8] ), .B(n314), .C(alu_op[2]), .D(
        n162), .Y(n1073) );
  AOI22X1 \myalu/muxs/m7/U3  ( .A(\myalu/s0[7] ), .B(n314), .C(alu_op[2]), .D(
        n161), .Y(n1072) );
  AOI22X1 \myalu/muxs/m6/U3  ( .A(\myalu/s0[6] ), .B(n314), .C(alu_op[2]), .D(
        n160), .Y(n1071) );
  AOI22X1 \myalu/muxs/m5/U3  ( .A(\myalu/s0[5] ), .B(n314), .C(alu_op[2]), .D(
        n159), .Y(n1070) );
  AOI22X1 \myalu/muxs/m4/U3  ( .A(\myalu/s0[4] ), .B(n314), .C(alu_op[2]), .D(
        n158), .Y(n1069) );
  AOI22X1 \myalu/muxs/m3/U3  ( .A(\myalu/s0[3] ), .B(n314), .C(alu_op[2]), .D(
        n157), .Y(n1068) );
  AOI22X1 \myalu/muxs/m2/U3  ( .A(\myalu/s0[2] ), .B(n314), .C(alu_op[2]), .D(
        n156), .Y(n1067) );
  AOI22X1 \myalu/muxs/m1/U3  ( .A(\myalu/s0[1] ), .B(n314), .C(alu_op[2]), .D(
        n155), .Y(n1066) );
  AOI22X1 \myalu/muxs/m0/U3  ( .A(\myalu/s0[0] ), .B(n314), .C(alu_op[2]), .D(
        n169), .Y(n1065) );
  AOI22X1 \myalu/mux0/m31/U3  ( .A(\myalu/s00[31] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[31] ), .Y(n1064) );
  AOI22X1 \myalu/mux0/m30/U3  ( .A(\myalu/s00[30] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[30] ), .Y(n1063) );
  AOI22X1 \myalu/mux0/m29/U3  ( .A(\myalu/s00[29] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[29] ), .Y(n1062) );
  AOI22X1 \myalu/mux0/m28/U3  ( .A(\myalu/s00[28] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[28] ), .Y(n1061) );
  AOI22X1 \myalu/mux0/m27/U3  ( .A(\myalu/s00[27] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[27] ), .Y(n1060) );
  AOI22X1 \myalu/mux0/m26/U3  ( .A(\myalu/s00[26] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[26] ), .Y(n1059) );
  AOI22X1 \myalu/mux0/m25/U3  ( .A(\myalu/s00[25] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[25] ), .Y(n1058) );
  AOI22X1 \myalu/mux0/m24/U3  ( .A(\myalu/s00[24] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[24] ), .Y(n1057) );
  AOI22X1 \myalu/mux0/m23/U3  ( .A(\myalu/s00[23] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[23] ), .Y(n1056) );
  AOI22X1 \myalu/mux0/m22/U3  ( .A(\myalu/s00[22] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[22] ), .Y(n1055) );
  AOI22X1 \myalu/mux0/m21/U3  ( .A(\myalu/s00[21] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[21] ), .Y(n1054) );
  AOI22X1 \myalu/mux0/m20/U3  ( .A(\myalu/s00[20] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[20] ), .Y(n1053) );
  AOI22X1 \myalu/mux0/m19/U3  ( .A(\myalu/s00[19] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[19] ), .Y(n1052) );
  AOI22X1 \myalu/mux0/m18/U3  ( .A(\myalu/s00[18] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[18] ), .Y(n1051) );
  AOI22X1 \myalu/mux0/m17/U3  ( .A(\myalu/s00[17] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[17] ), .Y(n1050) );
  AOI22X1 \myalu/mux0/m16/U3  ( .A(\myalu/s00[16] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[16] ), .Y(n1049) );
  AOI22X1 \myalu/mux0/m15/U3  ( .A(\myalu/s00[15] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[15] ), .Y(n1048) );
  AOI22X1 \myalu/mux0/m14/U3  ( .A(\myalu/s00[14] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[14] ), .Y(n1047) );
  AOI22X1 \myalu/mux0/m13/U3  ( .A(\myalu/s00[13] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[13] ), .Y(n1046) );
  AOI22X1 \myalu/mux0/m12/U3  ( .A(\myalu/s00[12] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[12] ), .Y(n1045) );
  AOI22X1 \myalu/mux0/m11/U3  ( .A(\myalu/s00[11] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[11] ), .Y(n1044) );
  AOI22X1 \myalu/mux0/m10/U3  ( .A(\myalu/s00[10] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[10] ), .Y(n1043) );
  AOI22X1 \myalu/mux0/m9/U3  ( .A(\myalu/s00[9] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[9] ), .Y(n1042) );
  AOI22X1 \myalu/mux0/m8/U3  ( .A(\myalu/s00[8] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[8] ), .Y(n1041) );
  AOI22X1 \myalu/mux0/m7/U3  ( .A(\myalu/s00[7] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[7] ), .Y(n1040) );
  AOI22X1 \myalu/mux0/m6/U3  ( .A(\myalu/s00[6] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[6] ), .Y(n1039) );
  AOI22X1 \myalu/mux0/m5/U3  ( .A(\myalu/s00[5] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[5] ), .Y(n1038) );
  AOI22X1 \myalu/mux0/m4/U3  ( .A(\myalu/s00[4] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[4] ), .Y(n1037) );
  AOI22X1 \myalu/mux0/m3/U3  ( .A(\myalu/s00[3] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[3] ), .Y(n1036) );
  AOI22X1 \myalu/mux0/m2/U3  ( .A(\myalu/s00[2] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[2] ), .Y(n1035) );
  AOI22X1 \myalu/mux0/m1/U3  ( .A(\myalu/s00[1] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[1] ), .Y(n1034) );
  AOI22X1 \myalu/mux0/m0/U3  ( .A(\myalu/s00[0] ), .B(n313), .C(alu_op[1]), 
        .D(\myalu/saddsub[0] ), .Y(n1033) );
  AOI22X1 \myalu/mux10/m31/U3  ( .A(\myalu/sand[31] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[31] ), .Y(n1032) );
  AOI22X1 \myalu/mux10/m30/U3  ( .A(\myalu/sand[30] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[30] ), .Y(n1031) );
  AOI22X1 \myalu/mux10/m29/U3  ( .A(\myalu/sand[29] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[29] ), .Y(n1030) );
  AOI22X1 \myalu/mux10/m28/U3  ( .A(\myalu/sand[28] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[28] ), .Y(n1029) );
  AOI22X1 \myalu/mux10/m27/U3  ( .A(\myalu/sand[27] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[27] ), .Y(n1028) );
  AOI22X1 \myalu/mux10/m26/U3  ( .A(\myalu/sand[26] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[26] ), .Y(n1027) );
  AOI22X1 \myalu/mux10/m25/U3  ( .A(\myalu/sand[25] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[25] ), .Y(n1026) );
  AOI22X1 \myalu/mux10/m24/U3  ( .A(\myalu/sand[24] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[24] ), .Y(n1025) );
  AOI22X1 \myalu/mux10/m23/U3  ( .A(\myalu/sand[23] ), .B(n312), .C(n310), .D(
        \myalu/sxnor[23] ), .Y(n1024) );
  AOI22X1 \myalu/mux10/m22/U3  ( .A(\myalu/sand[22] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[22] ), .Y(n1023) );
  AOI22X1 \myalu/mux10/m21/U3  ( .A(\myalu/sand[21] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[21] ), .Y(n1022) );
  AOI22X1 \myalu/mux10/m20/U3  ( .A(\myalu/sand[20] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[20] ), .Y(n1021) );
  AOI22X1 \myalu/mux10/m19/U3  ( .A(\myalu/sand[19] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[19] ), .Y(n1020) );
  AOI22X1 \myalu/mux10/m18/U3  ( .A(\myalu/sand[18] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[18] ), .Y(n1019) );
  AOI22X1 \myalu/mux10/m17/U3  ( .A(\myalu/sand[17] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[17] ), .Y(n1018) );
  AOI22X1 \myalu/mux10/m16/U3  ( .A(\myalu/sand[16] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[16] ), .Y(n1017) );
  AOI22X1 \myalu/mux10/m15/U3  ( .A(\myalu/sand[15] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[15] ), .Y(n1016) );
  AOI22X1 \myalu/mux10/m14/U3  ( .A(\myalu/sand[14] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[14] ), .Y(n1015) );
  AOI22X1 \myalu/mux10/m13/U3  ( .A(\myalu/sand[13] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[13] ), .Y(n1014) );
  AOI22X1 \myalu/mux10/m12/U3  ( .A(\myalu/sand[12] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[12] ), .Y(n1013) );
  AOI22X1 \myalu/mux10/m11/U3  ( .A(\myalu/sand[11] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[11] ), .Y(n1012) );
  AOI22X1 \myalu/mux10/m10/U3  ( .A(\myalu/sand[10] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[10] ), .Y(n1011) );
  AOI22X1 \myalu/mux10/m9/U3  ( .A(\myalu/sand[9] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[9] ), .Y(n1010) );
  AOI22X1 \myalu/mux10/m8/U3  ( .A(\myalu/sand[8] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[8] ), .Y(n1009) );
  AOI22X1 \myalu/mux10/m7/U3  ( .A(\myalu/sand[7] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[7] ), .Y(n1008) );
  AOI22X1 \myalu/mux10/m6/U3  ( .A(\myalu/sand[6] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[6] ), .Y(n1007) );
  AOI22X1 \myalu/mux10/m5/U3  ( .A(\myalu/sand[5] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[5] ), .Y(n1006) );
  AOI22X1 \myalu/mux10/m4/U3  ( .A(\myalu/sand[4] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[4] ), .Y(n1005) );
  AOI22X1 \myalu/mux10/m3/U3  ( .A(\myalu/sand[3] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[3] ), .Y(n1004) );
  AOI22X1 \myalu/mux10/m2/U3  ( .A(\myalu/sand[2] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[2] ), .Y(n1003) );
  AOI22X1 \myalu/mux10/m1/U3  ( .A(\myalu/sand[1] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[1] ), .Y(n1002) );
  AOI22X1 \myalu/mux10/m0/U3  ( .A(\myalu/sand[0] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/sxnor[0] ), .Y(n1001) );
  AOI22X1 \myalu/mux00/m31/U3  ( .A(\myalu/ssl[31] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[31] ), .Y(n1000) );
  AOI22X1 \myalu/mux00/m30/U3  ( .A(\myalu/ssl[30] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[30] ), .Y(n999) );
  AOI22X1 \myalu/mux00/m29/U3  ( .A(\myalu/ssl[29] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[29] ), .Y(n998) );
  AOI22X1 \myalu/mux00/m28/U3  ( .A(\myalu/ssl[28] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[28] ), .Y(n997) );
  AOI22X1 \myalu/mux00/m27/U3  ( .A(\myalu/ssl[27] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[27] ), .Y(n996) );
  AOI22X1 \myalu/mux00/m26/U3  ( .A(\myalu/ssl[26] ), .B(n312), .C(n310), .D(
        \myalu/ssr[26] ), .Y(n995) );
  AOI22X1 \myalu/mux00/m25/U3  ( .A(\myalu/ssl[25] ), .B(n312), .C(n309), .D(
        \myalu/ssr[25] ), .Y(n994) );
  AOI22X1 \myalu/mux00/m24/U3  ( .A(\myalu/ssl[24] ), .B(n312), .C(n308), .D(
        \myalu/ssr[24] ), .Y(n993) );
  AOI22X1 \myalu/mux00/m23/U3  ( .A(\myalu/ssl[23] ), .B(n312), .C(n309), .D(
        \myalu/ssr[23] ), .Y(n992) );
  AOI22X1 \myalu/mux00/m22/U3  ( .A(\myalu/ssl[22] ), .B(n312), .C(n308), .D(
        \myalu/ssr[22] ), .Y(n991) );
  AOI22X1 \myalu/mux00/m21/U3  ( .A(\myalu/ssl[21] ), .B(n312), .C(n309), .D(
        \myalu/ssr[21] ), .Y(n990) );
  AOI22X1 \myalu/mux00/m20/U3  ( .A(\myalu/ssl[20] ), .B(n312), .C(n308), .D(
        \myalu/ssr[20] ), .Y(n989) );
  AOI22X1 \myalu/mux00/m19/U3  ( .A(\myalu/ssl[19] ), .B(n312), .C(n309), .D(
        \myalu/ssr[19] ), .Y(n988) );
  AOI22X1 \myalu/mux00/m18/U3  ( .A(\myalu/ssl[18] ), .B(n312), .C(n308), .D(
        \myalu/ssr[18] ), .Y(n987) );
  AOI22X1 \myalu/mux00/m17/U3  ( .A(\myalu/ssl[17] ), .B(n312), .C(n309), .D(
        \myalu/ssr[17] ), .Y(n986) );
  AOI22X1 \myalu/mux00/m16/U3  ( .A(\myalu/ssl[16] ), .B(n312), .C(n308), .D(
        \myalu/ssr[16] ), .Y(n985) );
  AOI22X1 \myalu/mux00/m15/U3  ( .A(\myalu/ssl[15] ), .B(n312), .C(n309), .D(
        \myalu/ssr[15] ), .Y(n984) );
  AOI22X1 \myalu/mux00/m14/U3  ( .A(\myalu/ssl[14] ), .B(n312), .C(n308), .D(
        \myalu/ssr[14] ), .Y(n983) );
  AOI22X1 \myalu/mux00/m13/U3  ( .A(\myalu/ssl[13] ), .B(n312), .C(n309), .D(
        \myalu/ssr[13] ), .Y(n982) );
  AOI22X1 \myalu/mux00/m12/U3  ( .A(\myalu/ssl[12] ), .B(n312), .C(n308), .D(
        \myalu/ssr[12] ), .Y(n981) );
  AOI22X1 \myalu/mux00/m11/U3  ( .A(\myalu/ssl[11] ), .B(n312), .C(n309), .D(
        \myalu/ssr[11] ), .Y(n980) );
  AOI22X1 \myalu/mux00/m10/U3  ( .A(\myalu/ssl[10] ), .B(n312), .C(n308), .D(
        \myalu/ssr[10] ), .Y(n979) );
  AOI22X1 \myalu/mux00/m9/U3  ( .A(\myalu/ssl[9] ), .B(n312), .C(alu_op[0]), 
        .D(\myalu/ssr[9] ), .Y(n978) );
  AOI22X1 \myalu/mux00/m8/U3  ( .A(\myalu/ssl[8] ), .B(n312), .C(n308), .D(
        \myalu/ssr[8] ), .Y(n977) );
  AOI22X1 \myalu/mux00/m7/U3  ( .A(\myalu/ssl[7] ), .B(n312), .C(n308), .D(
        \myalu/ssr[7] ), .Y(n976) );
  AOI22X1 \myalu/mux00/m6/U3  ( .A(\myalu/ssl[6] ), .B(n312), .C(n308), .D(
        \myalu/ssr[6] ), .Y(n975) );
  AOI22X1 \myalu/mux00/m5/U3  ( .A(\myalu/ssl[5] ), .B(n312), .C(n308), .D(
        \myalu/ssr[5] ), .Y(n974) );
  AOI22X1 \myalu/mux00/m4/U3  ( .A(\myalu/ssl[4] ), .B(n312), .C(n308), .D(
        \myalu/ssr[4] ), .Y(n973) );
  AOI22X1 \myalu/mux00/m3/U3  ( .A(\myalu/ssl[3] ), .B(n312), .C(n308), .D(
        \myalu/ssr[3] ), .Y(n972) );
  AOI22X1 \myalu/mux00/m2/U3  ( .A(\myalu/ssl[2] ), .B(n312), .C(n308), .D(
        \myalu/ssr[2] ), .Y(n971) );
  AOI22X1 \myalu/mux00/m1/U3  ( .A(\myalu/ssl[1] ), .B(n312), .C(n310), .D(
        \myalu/ssr[1] ), .Y(n970) );
  AOI22X1 \myalu/mux00/m0/U3  ( .A(\myalu/ssl[0] ), .B(n311), .C(alu_op[0]), 
        .D(\myalu/ssr[0] ), .Y(n969) );
  AOI22X1 \mypc/mux1/m7/U3  ( .A(\mypc/temp_pc0[7] ), .B(n961), .C(n211), .D(
        pc[7]), .Y(n968) );
  AOI22X1 \mypc/mux1/m6/U3  ( .A(\mypc/temp_pc0[6] ), .B(n961), .C(n211), .D(
        pc[6]), .Y(n967) );
  AOI22X1 \mypc/mux1/m5/U3  ( .A(\mypc/temp_pc0[5] ), .B(n961), .C(n211), .D(
        pc[5]), .Y(n966) );
  AOI22X1 \mypc/mux1/m4/U3  ( .A(\mypc/temp_pc0[4] ), .B(n961), .C(n211), .D(
        pc[4]), .Y(n965) );
  AOI22X1 \mypc/mux1/m3/U3  ( .A(\mypc/temp_pc0[3] ), .B(n961), .C(n211), .D(
        pc[3]), .Y(n964) );
  AOI22X1 \mypc/mux1/m2/U3  ( .A(\mypc/temp_pc0[2] ), .B(n961), .C(n211), .D(
        pc[2]), .Y(n963) );
  AOI22X1 \mypc/mux1/m1/U3  ( .A(\mypc/temp_pc0[1] ), .B(n961), .C(n211), .D(
        pc[1]), .Y(n962) );
  AOI22X1 \mypc/mux1/m0/U3  ( .A(\mypc/temp_pc0[0] ), .B(n961), .C(n211), .D(
        pc[0]), .Y(n960) );
  AOI22X1 \mypc/mux0/m7/U3  ( .A(\mypc/inc_pc[7] ), .B(n952), .C(
        \mypc/branch_en ), .D(addr_s[3]), .Y(n959) );
  AOI22X1 \mypc/mux0/m6/U3  ( .A(\mypc/inc_pc[6] ), .B(n952), .C(
        \mypc/branch_en ), .D(addr_s[2]), .Y(n958) );
  AOI22X1 \mypc/mux0/m5/U3  ( .A(\mypc/inc_pc[5] ), .B(n952), .C(
        \mypc/branch_en ), .D(n210), .Y(n957) );
  AOI22X1 \mypc/mux0/m4/U3  ( .A(\mypc/inc_pc[4] ), .B(n952), .C(
        \mypc/branch_en ), .D(n209), .Y(n956) );
  AOI22X1 \mypc/mux0/m3/U3  ( .A(\mypc/inc_pc[3] ), .B(n952), .C(
        \mypc/branch_en ), .D(\myram/db/en1 ), .Y(n955) );
  AOI22X1 \mypc/mux0/m2/U3  ( .A(\mypc/inc_pc[2] ), .B(n952), .C(
        \mypc/branch_en ), .D(addr_b[2]), .Y(n954) );
  AOI22X1 \mypc/mux0/m1/U3  ( .A(\mypc/inc_pc[1] ), .B(n952), .C(
        \mypc/branch_en ), .D(n206), .Y(n953) );
  AOI22X1 \mypc/mux0/m0/U3  ( .A(\mypc/inc_pc[0] ), .B(n952), .C(
        \mypc/branch_en ), .D(n205), .Y(n951) );
  AOI22X1 \alu_out/m7/U3  ( .A(alu_s[7]), .B(n315), .C(imm_en), .D(
        \myram/da/en1 ), .Y(n949) );
  AOI22X1 \alu_out/m6/U3  ( .A(alu_s[6]), .B(n315), .C(imm_en), .D(addr_a[2]), 
        .Y(n948) );
  AOI22X1 \alu_out/m5/U3  ( .A(alu_s[5]), .B(n315), .C(imm_en), .D(n208), .Y(
        n947) );
  AOI22X1 \alu_out/m4/U3  ( .A(alu_s[4]), .B(n315), .C(imm_en), .D(n207), .Y(
        n946) );
  AOI22X1 \alu_out/m3/U3  ( .A(alu_s[3]), .B(n315), .C(imm_en), .D(
        \myram/db/en1 ), .Y(n945) );
  AOI22X1 \alu_out/m2/U3  ( .A(alu_s[2]), .B(n315), .C(imm_en), .D(addr_b[2]), 
        .Y(n944) );
  AOI22X1 \alu_out/m1/U3  ( .A(alu_s[1]), .B(n315), .C(imm_en), .D(n206), .Y(
        n943) );
  DFFPOSX1 \myram/m0/d/d31/q_reg  ( .D(\myram/m0/mux_out[31] ), .CLK(clk), .Q(
        \myram/m0/dout[31] ) );
  DFFPOSX1 \myram/m0/d/d30/q_reg  ( .D(\myram/m0/mux_out[30] ), .CLK(clk), .Q(
        \myram/m0/dout[30] ) );
  DFFPOSX1 \myram/m0/d/d29/q_reg  ( .D(\myram/m0/mux_out[29] ), .CLK(clk), .Q(
        \myram/m0/dout[29] ) );
  DFFPOSX1 \myram/m0/d/d28/q_reg  ( .D(\myram/m0/mux_out[28] ), .CLK(clk), .Q(
        \myram/m0/dout[28] ) );
  DFFPOSX1 \myram/m0/d/d27/q_reg  ( .D(\myram/m0/mux_out[27] ), .CLK(clk), .Q(
        \myram/m0/dout[27] ) );
  DFFPOSX1 \myram/m0/d/d26/q_reg  ( .D(\myram/m0/mux_out[26] ), .CLK(clk), .Q(
        \myram/m0/dout[26] ) );
  DFFPOSX1 \myram/m0/d/d25/q_reg  ( .D(\myram/m0/mux_out[25] ), .CLK(clk), .Q(
        \myram/m0/dout[25] ) );
  DFFPOSX1 \myram/m0/d/d24/q_reg  ( .D(\myram/m0/mux_out[24] ), .CLK(clk), .Q(
        \myram/m0/dout[24] ) );
  DFFPOSX1 \myram/m0/d/d23/q_reg  ( .D(\myram/m0/mux_out[23] ), .CLK(clk), .Q(
        \myram/m0/dout[23] ) );
  DFFPOSX1 \myram/m0/d/d22/q_reg  ( .D(\myram/m0/mux_out[22] ), .CLK(clk), .Q(
        \myram/m0/dout[22] ) );
  DFFPOSX1 \myram/m0/d/d21/q_reg  ( .D(\myram/m0/mux_out[21] ), .CLK(clk), .Q(
        \myram/m0/dout[21] ) );
  DFFPOSX1 \myram/m0/d/d20/q_reg  ( .D(\myram/m0/mux_out[20] ), .CLK(clk), .Q(
        \myram/m0/dout[20] ) );
  DFFPOSX1 \myram/m0/d/d19/q_reg  ( .D(\myram/m0/mux_out[19] ), .CLK(clk), .Q(
        \myram/m0/dout[19] ) );
  DFFPOSX1 \myram/m0/d/d18/q_reg  ( .D(\myram/m0/mux_out[18] ), .CLK(clk), .Q(
        \myram/m0/dout[18] ) );
  DFFPOSX1 \myram/m0/d/d17/q_reg  ( .D(\myram/m0/mux_out[17] ), .CLK(clk), .Q(
        \myram/m0/dout[17] ) );
  DFFPOSX1 \myram/m0/d/d16/q_reg  ( .D(\myram/m0/mux_out[16] ), .CLK(clk), .Q(
        \myram/m0/dout[16] ) );
  DFFPOSX1 \myram/m0/d/d15/q_reg  ( .D(\myram/m0/mux_out[15] ), .CLK(clk), .Q(
        \myram/m0/dout[15] ) );
  DFFPOSX1 \myram/m0/d/d14/q_reg  ( .D(\myram/m0/mux_out[14] ), .CLK(clk), .Q(
        \myram/m0/dout[14] ) );
  DFFPOSX1 \myram/m0/d/d13/q_reg  ( .D(\myram/m0/mux_out[13] ), .CLK(clk), .Q(
        \myram/m0/dout[13] ) );
  DFFPOSX1 \myram/m0/d/d12/q_reg  ( .D(\myram/m0/mux_out[12] ), .CLK(clk), .Q(
        \myram/m0/dout[12] ) );
  DFFPOSX1 \myram/m0/d/d11/q_reg  ( .D(\myram/m0/mux_out[11] ), .CLK(clk), .Q(
        \myram/m0/dout[11] ) );
  DFFPOSX1 \myram/m0/d/d10/q_reg  ( .D(\myram/m0/mux_out[10] ), .CLK(clk), .Q(
        \myram/m0/dout[10] ) );
  DFFPOSX1 \myram/m0/d/d9/q_reg  ( .D(\myram/m0/mux_out[9] ), .CLK(clk), .Q(
        \myram/m0/dout[9] ) );
  DFFPOSX1 \myram/m0/d/d8/q_reg  ( .D(\myram/m0/mux_out[8] ), .CLK(clk), .Q(
        \myram/m0/dout[8] ) );
  DFFPOSX1 \myram/m0/d/d7/q_reg  ( .D(\myram/m0/mux_out[7] ), .CLK(clk), .Q(
        \myram/m0/dout[7] ) );
  DFFPOSX1 \myram/m0/d/d6/q_reg  ( .D(\myram/m0/mux_out[6] ), .CLK(clk), .Q(
        \myram/m0/dout[6] ) );
  DFFPOSX1 \myram/m0/d/d5/q_reg  ( .D(\myram/m0/mux_out[5] ), .CLK(clk), .Q(
        \myram/m0/dout[5] ) );
  DFFPOSX1 \myram/m0/d/d4/q_reg  ( .D(\myram/m0/mux_out[4] ), .CLK(clk), .Q(
        \myram/m0/dout[4] ) );
  DFFPOSX1 \myram/m0/d/d3/q_reg  ( .D(\myram/m0/mux_out[3] ), .CLK(clk), .Q(
        \myram/m0/dout[3] ) );
  DFFPOSX1 \myram/m0/d/d2/q_reg  ( .D(\myram/m0/mux_out[2] ), .CLK(clk), .Q(
        \myram/m0/dout[2] ) );
  DFFPOSX1 \myram/m0/d/d1/q_reg  ( .D(\myram/m0/mux_out[1] ), .CLK(clk), .Q(
        \myram/m0/dout[1] ) );
  DFFPOSX1 \myram/m0/d/d0/q_reg  ( .D(\myram/m0/mux_out[0] ), .CLK(clk), .Q(
        \myram/m0/dout[0] ) );
  DFFPOSX1 \mypc/d/d7/q_reg  ( .D(next_pc[7]), .CLK(clk), .Q(pc[7]) );
  DFFPOSX1 \mypc/d/d6/q_reg  ( .D(next_pc[6]), .CLK(clk), .Q(pc[6]) );
  DFFPOSX1 \mypc/d/d5/q_reg  ( .D(next_pc[5]), .CLK(clk), .Q(pc[5]) );
  DFFPOSX1 \mypc/d/d4/q_reg  ( .D(next_pc[4]), .CLK(clk), .Q(pc[4]) );
  DFFPOSX1 \mypc/d/d3/q_reg  ( .D(next_pc[3]), .CLK(clk), .Q(pc[3]) );
  DFFPOSX1 \mypc/d/d2/q_reg  ( .D(next_pc[2]), .CLK(clk), .Q(pc[2]) );
  DFFPOSX1 \mypc/d/d1/q_reg  ( .D(next_pc[1]), .CLK(clk), .Q(pc[1]) );
  XNOR2X1 \myalu/myadder/myadder/a31/U5  ( .A(a[31]), .B(
        \myalu/myadder/xb[31] ), .Y(n942) );
  XOR2X1 \myalu/myadder/myadder/a31/U2  ( .A(n941), .B(n942), .Y(
        \myalu/saddsub[31] ) );
  XNOR2X1 \myalu/myadder/myadder/a30/U5  ( .A(a[30]), .B(
        \myalu/myadder/xb[30] ), .Y(n939) );
  OAI21X1 \myalu/myadder/myadder/a30/U3  ( .A(n939), .B(n938), .C(n120), .Y(
        \myalu/myadder/myadder/c31 ) );
  XOR2X1 \myalu/myadder/myadder/a30/U2  ( .A(n938), .B(n939), .Y(
        \myalu/saddsub[30] ) );
  XNOR2X1 \myalu/myadder/myadder/a29/U5  ( .A(a[29]), .B(
        \myalu/myadder/xb[29] ), .Y(n936) );
  OAI21X1 \myalu/myadder/myadder/a29/U3  ( .A(n936), .B(n935), .C(n91), .Y(
        \myalu/myadder/myadder/c30 ) );
  XOR2X1 \myalu/myadder/myadder/a29/U2  ( .A(n935), .B(n936), .Y(
        \myalu/saddsub[29] ) );
  XNOR2X1 \myalu/myadder/myadder/a28/U5  ( .A(a[28]), .B(
        \myalu/myadder/xb[28] ), .Y(n933) );
  OAI21X1 \myalu/myadder/myadder/a28/U3  ( .A(n933), .B(n932), .C(n79), .Y(
        \myalu/myadder/myadder/c29 ) );
  XOR2X1 \myalu/myadder/myadder/a28/U2  ( .A(n932), .B(n933), .Y(
        \myalu/saddsub[28] ) );
  XNOR2X1 \myalu/myadder/myadder/a27/U5  ( .A(a[27]), .B(
        \myalu/myadder/xb[27] ), .Y(n930) );
  OAI21X1 \myalu/myadder/myadder/a27/U3  ( .A(n930), .B(n929), .C(n118), .Y(
        \myalu/myadder/myadder/c28 ) );
  XOR2X1 \myalu/myadder/myadder/a27/U2  ( .A(n929), .B(n930), .Y(
        \myalu/saddsub[27] ) );
  XNOR2X1 \myalu/myadder/myadder/a26/U5  ( .A(a[26]), .B(
        \myalu/myadder/xb[26] ), .Y(n927) );
  OAI21X1 \myalu/myadder/myadder/a26/U3  ( .A(n927), .B(n926), .C(n102), .Y(
        \myalu/myadder/myadder/c27 ) );
  XOR2X1 \myalu/myadder/myadder/a26/U2  ( .A(n926), .B(n927), .Y(
        \myalu/saddsub[26] ) );
  XNOR2X1 \myalu/myadder/myadder/a25/U5  ( .A(a[25]), .B(
        \myalu/myadder/xb[25] ), .Y(n924) );
  OAI21X1 \myalu/myadder/myadder/a25/U3  ( .A(n924), .B(n923), .C(n89), .Y(
        \myalu/myadder/myadder/c26 ) );
  XOR2X1 \myalu/myadder/myadder/a25/U2  ( .A(n923), .B(n924), .Y(
        \myalu/saddsub[25] ) );
  XNOR2X1 \myalu/myadder/myadder/a24/U5  ( .A(a[24]), .B(
        \myalu/myadder/xb[24] ), .Y(n921) );
  OAI21X1 \myalu/myadder/myadder/a24/U3  ( .A(n921), .B(n920), .C(n116), .Y(
        \myalu/myadder/myadder/c25 ) );
  XOR2X1 \myalu/myadder/myadder/a24/U2  ( .A(n920), .B(n921), .Y(
        \myalu/saddsub[24] ) );
  XNOR2X1 \myalu/myadder/myadder/a23/U5  ( .A(a[23]), .B(
        \myalu/myadder/xb[23] ), .Y(n918) );
  OAI21X1 \myalu/myadder/myadder/a23/U3  ( .A(n918), .B(n917), .C(n101), .Y(
        \myalu/myadder/myadder/c24 ) );
  XOR2X1 \myalu/myadder/myadder/a23/U2  ( .A(n917), .B(n918), .Y(
        \myalu/saddsub[23] ) );
  XNOR2X1 \myalu/myadder/myadder/a22/U5  ( .A(a[22]), .B(
        \myalu/myadder/xb[22] ), .Y(n915) );
  OAI21X1 \myalu/myadder/myadder/a22/U3  ( .A(n915), .B(n914), .C(n78), .Y(
        \myalu/myadder/myadder/c23 ) );
  XOR2X1 \myalu/myadder/myadder/a22/U2  ( .A(n914), .B(n915), .Y(
        \myalu/saddsub[22] ) );
  XNOR2X1 \myalu/myadder/myadder/a21/U5  ( .A(a[21]), .B(
        \myalu/myadder/xb[21] ), .Y(n912) );
  OAI21X1 \myalu/myadder/myadder/a21/U3  ( .A(n912), .B(n911), .C(n84), .Y(
        \myalu/myadder/myadder/c22 ) );
  XOR2X1 \myalu/myadder/myadder/a21/U2  ( .A(n911), .B(n912), .Y(
        \myalu/saddsub[21] ) );
  XNOR2X1 \myalu/myadder/myadder/a20/U5  ( .A(a[20]), .B(
        \myalu/myadder/xb[20] ), .Y(n909) );
  OAI21X1 \myalu/myadder/myadder/a20/U3  ( .A(n909), .B(n908), .C(n111), .Y(
        \myalu/myadder/myadder/c21 ) );
  XOR2X1 \myalu/myadder/myadder/a20/U2  ( .A(n908), .B(n909), .Y(
        \myalu/saddsub[20] ) );
  XNOR2X1 \myalu/myadder/myadder/a19/U5  ( .A(a[19]), .B(
        \myalu/myadder/xb[19] ), .Y(n906) );
  OAI21X1 \myalu/myadder/myadder/a19/U3  ( .A(n906), .B(n905), .C(n97), .Y(
        \myalu/myadder/myadder/c20 ) );
  XOR2X1 \myalu/myadder/myadder/a19/U2  ( .A(n905), .B(n906), .Y(
        \myalu/saddsub[19] ) );
  XNOR2X1 \myalu/myadder/myadder/a18/U5  ( .A(a[18]), .B(
        \myalu/myadder/xb[18] ), .Y(n903) );
  OAI21X1 \myalu/myadder/myadder/a18/U3  ( .A(n903), .B(n902), .C(n85), .Y(
        \myalu/myadder/myadder/c19 ) );
  XOR2X1 \myalu/myadder/myadder/a18/U2  ( .A(n902), .B(n903), .Y(
        \myalu/saddsub[18] ) );
  XNOR2X1 \myalu/myadder/myadder/a17/U5  ( .A(a[17]), .B(
        \myalu/myadder/xb[17] ), .Y(n900) );
  OAI21X1 \myalu/myadder/myadder/a17/U3  ( .A(n900), .B(n899), .C(n112), .Y(
        \myalu/myadder/myadder/c18 ) );
  XOR2X1 \myalu/myadder/myadder/a17/U2  ( .A(n899), .B(n900), .Y(
        \myalu/saddsub[17] ) );
  XNOR2X1 \myalu/myadder/myadder/a16/U5  ( .A(a[16]), .B(
        \myalu/myadder/xb[16] ), .Y(n897) );
  OAI21X1 \myalu/myadder/myadder/a16/U3  ( .A(n897), .B(n896), .C(n98), .Y(
        \myalu/myadder/myadder/c17 ) );
  XOR2X1 \myalu/myadder/myadder/a16/U2  ( .A(n896), .B(n897), .Y(
        \myalu/saddsub[16] ) );
  XNOR2X1 \myalu/myadder/myadder/a15/U5  ( .A(a[15]), .B(
        \myalu/myadder/xb[15] ), .Y(n894) );
  OAI21X1 \myalu/myadder/myadder/a15/U3  ( .A(n894), .B(n893), .C(n86), .Y(
        \myalu/myadder/myadder/c16 ) );
  XOR2X1 \myalu/myadder/myadder/a15/U2  ( .A(n893), .B(n894), .Y(
        \myalu/saddsub[15] ) );
  XNOR2X1 \myalu/myadder/myadder/a14/U5  ( .A(a[14]), .B(
        \myalu/myadder/xb[14] ), .Y(n891) );
  OAI21X1 \myalu/myadder/myadder/a14/U3  ( .A(n891), .B(n890), .C(n113), .Y(
        \myalu/myadder/myadder/c15 ) );
  XOR2X1 \myalu/myadder/myadder/a14/U2  ( .A(n890), .B(n891), .Y(
        \myalu/saddsub[14] ) );
  XNOR2X1 \myalu/myadder/myadder/a13/U5  ( .A(a[13]), .B(
        \myalu/myadder/xb[13] ), .Y(n888) );
  OAI21X1 \myalu/myadder/myadder/a13/U3  ( .A(n888), .B(n887), .C(n99), .Y(
        \myalu/myadder/myadder/c14 ) );
  XOR2X1 \myalu/myadder/myadder/a13/U2  ( .A(n887), .B(n888), .Y(
        \myalu/saddsub[13] ) );
  XNOR2X1 \myalu/myadder/myadder/a12/U5  ( .A(a[12]), .B(
        \myalu/myadder/xb[12] ), .Y(n885) );
  OAI21X1 \myalu/myadder/myadder/a12/U3  ( .A(n885), .B(n884), .C(n87), .Y(
        \myalu/myadder/myadder/c13 ) );
  XOR2X1 \myalu/myadder/myadder/a12/U2  ( .A(n884), .B(n885), .Y(
        \myalu/saddsub[12] ) );
  XNOR2X1 \myalu/myadder/myadder/a11/U5  ( .A(a[11]), .B(
        \myalu/myadder/xb[11] ), .Y(n882) );
  OAI21X1 \myalu/myadder/myadder/a11/U3  ( .A(n882), .B(n881), .C(n114), .Y(
        \myalu/myadder/myadder/c12 ) );
  XOR2X1 \myalu/myadder/myadder/a11/U2  ( .A(n881), .B(n882), .Y(
        \myalu/saddsub[11] ) );
  XNOR2X1 \myalu/myadder/myadder/a10/U5  ( .A(a[10]), .B(
        \myalu/myadder/xb[10] ), .Y(n879) );
  OAI21X1 \myalu/myadder/myadder/a10/U3  ( .A(n879), .B(n878), .C(n100), .Y(
        \myalu/myadder/myadder/c11 ) );
  XOR2X1 \myalu/myadder/myadder/a10/U2  ( .A(n878), .B(n879), .Y(
        \myalu/saddsub[10] ) );
  XNOR2X1 \myalu/myadder/myadder/a9/U5  ( .A(a[9]), .B(\myalu/myadder/xb[9] ), 
        .Y(n876) );
  OAI21X1 \myalu/myadder/myadder/a9/U3  ( .A(n876), .B(n875), .C(n88), .Y(
        \myalu/myadder/myadder/c10 ) );
  XOR2X1 \myalu/myadder/myadder/a9/U2  ( .A(n875), .B(n876), .Y(
        \myalu/saddsub[9] ) );
  XNOR2X1 \myalu/myadder/myadder/a8/U5  ( .A(a[8]), .B(\myalu/myadder/xb[8] ), 
        .Y(n873) );
  OAI21X1 \myalu/myadder/myadder/a8/U3  ( .A(n873), .B(n872), .C(n119), .Y(
        \myalu/myadder/myadder/c9 ) );
  XOR2X1 \myalu/myadder/myadder/a8/U2  ( .A(n872), .B(n873), .Y(
        \myalu/saddsub[8] ) );
  XNOR2X1 \myalu/myadder/myadder/a7/U5  ( .A(a[7]), .B(\myalu/myadder/xb[7] ), 
        .Y(n870) );
  OAI21X1 \myalu/myadder/myadder/a7/U3  ( .A(n870), .B(n869), .C(n103), .Y(
        \myalu/myadder/myadder/c8 ) );
  XOR2X1 \myalu/myadder/myadder/a7/U2  ( .A(n869), .B(n870), .Y(
        \myalu/saddsub[7] ) );
  XNOR2X1 \myalu/myadder/myadder/a6/U5  ( .A(a[6]), .B(\myalu/myadder/xb[6] ), 
        .Y(n867) );
  OAI21X1 \myalu/myadder/myadder/a6/U3  ( .A(n867), .B(n866), .C(n90), .Y(
        \myalu/myadder/myadder/c7 ) );
  XOR2X1 \myalu/myadder/myadder/a6/U2  ( .A(n866), .B(n867), .Y(
        \myalu/saddsub[6] ) );
  XNOR2X1 \myalu/myadder/myadder/a5/U5  ( .A(a[5]), .B(\myalu/myadder/xb[5] ), 
        .Y(n864) );
  OAI21X1 \myalu/myadder/myadder/a5/U3  ( .A(n864), .B(n863), .C(n115), .Y(
        \myalu/myadder/myadder/c6 ) );
  XOR2X1 \myalu/myadder/myadder/a5/U2  ( .A(n863), .B(n864), .Y(
        \myalu/saddsub[5] ) );
  XNOR2X1 \myalu/myadder/myadder/a4/U5  ( .A(a[4]), .B(\myalu/myadder/xb[4] ), 
        .Y(n861) );
  OAI21X1 \myalu/myadder/myadder/a4/U3  ( .A(n861), .B(n860), .C(n95), .Y(
        \myalu/myadder/myadder/c5 ) );
  XOR2X1 \myalu/myadder/myadder/a4/U2  ( .A(n860), .B(n861), .Y(
        \myalu/saddsub[4] ) );
  XNOR2X1 \myalu/myadder/myadder/a3/U5  ( .A(a[3]), .B(\myalu/myadder/xb[3] ), 
        .Y(n858) );
  OAI21X1 \myalu/myadder/myadder/a3/U3  ( .A(n858), .B(n857), .C(n77), .Y(
        \myalu/myadder/myadder/c4 ) );
  XOR2X1 \myalu/myadder/myadder/a3/U2  ( .A(n857), .B(n858), .Y(
        \myalu/saddsub[3] ) );
  XNOR2X1 \myalu/myadder/myadder/a2/U5  ( .A(a[2]), .B(\myalu/myadder/xb[2] ), 
        .Y(n855) );
  OAI21X1 \myalu/myadder/myadder/a2/U3  ( .A(n855), .B(n854), .C(n83), .Y(
        \myalu/myadder/myadder/c3 ) );
  XOR2X1 \myalu/myadder/myadder/a2/U2  ( .A(n854), .B(n855), .Y(
        \myalu/saddsub[2] ) );
  XNOR2X1 \myalu/myadder/myadder/a1/U5  ( .A(a[1]), .B(\myalu/myadder/xb[1] ), 
        .Y(n852) );
  OAI21X1 \myalu/myadder/myadder/a1/U3  ( .A(n852), .B(n851), .C(n96), .Y(
        \myalu/myadder/myadder/c2 ) );
  XOR2X1 \myalu/myadder/myadder/a1/U2  ( .A(n851), .B(n852), .Y(
        \myalu/saddsub[1] ) );
  XNOR2X1 \myalu/myadder/myadder/a0/U5  ( .A(a[0]), .B(\myalu/myadder/xb[0] ), 
        .Y(n849) );
  OAI21X1 \myalu/myadder/myadder/a0/U3  ( .A(n849), .B(n311), .C(n117), .Y(
        \myalu/myadder/myadder/c1 ) );
  XOR2X1 \myalu/myadder/myadder/a0/U2  ( .A(n312), .B(n849), .Y(
        \myalu/saddsub[0] ) );
  XOR2X1 \mypc/myinc/a7/U2  ( .A(n190), .B(n848), .Y(\mypc/inc_pc[7] ) );
  XOR2X1 \mypc/myinc/a6/U2  ( .A(n189), .B(n847), .Y(\mypc/inc_pc[6] ) );
  XOR2X1 \mypc/myinc/a5/U2  ( .A(n188), .B(n846), .Y(\mypc/inc_pc[5] ) );
  XOR2X1 \mypc/myinc/a4/U2  ( .A(n187), .B(n845), .Y(\mypc/inc_pc[4] ) );
  XOR2X1 \mypc/myinc/a3/U2  ( .A(n184), .B(n844), .Y(\mypc/inc_pc[3] ) );
  XOR2X1 \mypc/myinc/a2/U2  ( .A(n186), .B(n843), .Y(\mypc/inc_pc[2] ) );
  XOR2X1 \mypc/myinc/a1/U2  ( .A(\mypc/inc_pc[0] ), .B(n842), .Y(
        \mypc/inc_pc[1] ) );
  DFFPOSX1 \myram/m15/d/d0/q_reg  ( .D(\myram/m15/mux_out[0] ), .CLK(clk), .Q(
        \myram/m15/dout[0] ) );
  DFFPOSX1 \myram/m15/d/d1/q_reg  ( .D(\myram/m15/mux_out[1] ), .CLK(clk), .Q(
        \myram/m15/dout[1] ) );
  DFFPOSX1 \myram/m15/d/d2/q_reg  ( .D(\myram/m15/mux_out[2] ), .CLK(clk), .Q(
        \myram/m15/dout[2] ) );
  DFFPOSX1 \myram/m15/d/d3/q_reg  ( .D(\myram/m15/mux_out[3] ), .CLK(clk), .Q(
        \myram/m15/dout[3] ) );
  DFFPOSX1 \myram/m15/d/d4/q_reg  ( .D(\myram/m15/mux_out[4] ), .CLK(clk), .Q(
        \myram/m15/dout[4] ) );
  DFFPOSX1 \myram/m15/d/d5/q_reg  ( .D(\myram/m15/mux_out[5] ), .CLK(clk), .Q(
        \myram/m15/dout[5] ) );
  DFFPOSX1 \myram/m15/d/d6/q_reg  ( .D(\myram/m15/mux_out[6] ), .CLK(clk), .Q(
        \myram/m15/dout[6] ) );
  DFFPOSX1 \myram/m15/d/d7/q_reg  ( .D(\myram/m15/mux_out[7] ), .CLK(clk), .Q(
        \myram/m15/dout[7] ) );
  DFFPOSX1 \myram/m15/d/d8/q_reg  ( .D(\myram/m15/mux_out[8] ), .CLK(clk), .Q(
        \myram/m15/dout[8] ) );
  DFFPOSX1 \myram/m15/d/d9/q_reg  ( .D(\myram/m15/mux_out[9] ), .CLK(clk), .Q(
        \myram/m15/dout[9] ) );
  DFFPOSX1 \myram/m15/d/d10/q_reg  ( .D(\myram/m15/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m15/dout[10] ) );
  DFFPOSX1 \myram/m15/d/d11/q_reg  ( .D(\myram/m15/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m15/dout[11] ) );
  DFFPOSX1 \myram/m15/d/d12/q_reg  ( .D(\myram/m15/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m15/dout[12] ) );
  DFFPOSX1 \myram/m15/d/d13/q_reg  ( .D(\myram/m15/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m15/dout[13] ) );
  DFFPOSX1 \myram/m15/d/d14/q_reg  ( .D(\myram/m15/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m15/dout[14] ) );
  DFFPOSX1 \myram/m15/d/d15/q_reg  ( .D(\myram/m15/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m15/dout[15] ) );
  DFFPOSX1 \myram/m15/d/d16/q_reg  ( .D(\myram/m15/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m15/dout[16] ) );
  DFFPOSX1 \myram/m15/d/d17/q_reg  ( .D(\myram/m15/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m15/dout[17] ) );
  DFFPOSX1 \myram/m15/d/d18/q_reg  ( .D(\myram/m15/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m15/dout[18] ) );
  DFFPOSX1 \myram/m15/d/d19/q_reg  ( .D(\myram/m15/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m15/dout[19] ) );
  DFFPOSX1 \myram/m15/d/d20/q_reg  ( .D(\myram/m15/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m15/dout[20] ) );
  DFFPOSX1 \myram/m15/d/d21/q_reg  ( .D(\myram/m15/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m15/dout[21] ) );
  DFFPOSX1 \myram/m15/d/d22/q_reg  ( .D(\myram/m15/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m15/dout[22] ) );
  DFFPOSX1 \myram/m15/d/d23/q_reg  ( .D(\myram/m15/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m15/dout[23] ) );
  DFFPOSX1 \myram/m15/d/d24/q_reg  ( .D(\myram/m15/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m15/dout[24] ) );
  DFFPOSX1 \myram/m15/d/d25/q_reg  ( .D(\myram/m15/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m15/dout[25] ) );
  DFFPOSX1 \myram/m15/d/d26/q_reg  ( .D(\myram/m15/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m15/dout[26] ) );
  DFFPOSX1 \myram/m15/d/d27/q_reg  ( .D(\myram/m15/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m15/dout[27] ) );
  DFFPOSX1 \myram/m15/d/d28/q_reg  ( .D(\myram/m15/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m15/dout[28] ) );
  DFFPOSX1 \myram/m15/d/d29/q_reg  ( .D(\myram/m15/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m15/dout[29] ) );
  DFFPOSX1 \myram/m15/d/d30/q_reg  ( .D(\myram/m15/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m15/dout[30] ) );
  DFFPOSX1 \myram/m15/d/d31/q_reg  ( .D(\myram/m15/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m15/dout[31] ) );
  DFFPOSX1 \myram/m14/d/d0/q_reg  ( .D(\myram/m14/mux_out[0] ), .CLK(clk), .Q(
        \myram/m14/dout[0] ) );
  DFFPOSX1 \myram/m14/d/d1/q_reg  ( .D(\myram/m14/mux_out[1] ), .CLK(clk), .Q(
        \myram/m14/dout[1] ) );
  DFFPOSX1 \myram/m14/d/d2/q_reg  ( .D(\myram/m14/mux_out[2] ), .CLK(clk), .Q(
        \myram/m14/dout[2] ) );
  DFFPOSX1 \myram/m14/d/d3/q_reg  ( .D(\myram/m14/mux_out[3] ), .CLK(clk), .Q(
        \myram/m14/dout[3] ) );
  DFFPOSX1 \myram/m14/d/d4/q_reg  ( .D(\myram/m14/mux_out[4] ), .CLK(clk), .Q(
        \myram/m14/dout[4] ) );
  DFFPOSX1 \myram/m14/d/d5/q_reg  ( .D(\myram/m14/mux_out[5] ), .CLK(clk), .Q(
        \myram/m14/dout[5] ) );
  DFFPOSX1 \myram/m14/d/d6/q_reg  ( .D(\myram/m14/mux_out[6] ), .CLK(clk), .Q(
        \myram/m14/dout[6] ) );
  DFFPOSX1 \myram/m14/d/d7/q_reg  ( .D(\myram/m14/mux_out[7] ), .CLK(clk), .Q(
        \myram/m14/dout[7] ) );
  DFFPOSX1 \myram/m14/d/d8/q_reg  ( .D(\myram/m14/mux_out[8] ), .CLK(clk), .Q(
        \myram/m14/dout[8] ) );
  DFFPOSX1 \myram/m14/d/d9/q_reg  ( .D(\myram/m14/mux_out[9] ), .CLK(clk), .Q(
        \myram/m14/dout[9] ) );
  DFFPOSX1 \myram/m14/d/d10/q_reg  ( .D(\myram/m14/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m14/dout[10] ) );
  DFFPOSX1 \myram/m14/d/d11/q_reg  ( .D(\myram/m14/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m14/dout[11] ) );
  DFFPOSX1 \myram/m14/d/d12/q_reg  ( .D(\myram/m14/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m14/dout[12] ) );
  DFFPOSX1 \myram/m14/d/d13/q_reg  ( .D(\myram/m14/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m14/dout[13] ) );
  DFFPOSX1 \myram/m14/d/d14/q_reg  ( .D(\myram/m14/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m14/dout[14] ) );
  DFFPOSX1 \myram/m14/d/d15/q_reg  ( .D(\myram/m14/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m14/dout[15] ) );
  DFFPOSX1 \myram/m14/d/d16/q_reg  ( .D(\myram/m14/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m14/dout[16] ) );
  DFFPOSX1 \myram/m14/d/d17/q_reg  ( .D(\myram/m14/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m14/dout[17] ) );
  DFFPOSX1 \myram/m14/d/d18/q_reg  ( .D(\myram/m14/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m14/dout[18] ) );
  DFFPOSX1 \myram/m14/d/d19/q_reg  ( .D(\myram/m14/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m14/dout[19] ) );
  DFFPOSX1 \myram/m14/d/d20/q_reg  ( .D(\myram/m14/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m14/dout[20] ) );
  DFFPOSX1 \myram/m14/d/d21/q_reg  ( .D(\myram/m14/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m14/dout[21] ) );
  DFFPOSX1 \myram/m14/d/d22/q_reg  ( .D(\myram/m14/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m14/dout[22] ) );
  DFFPOSX1 \myram/m14/d/d23/q_reg  ( .D(\myram/m14/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m14/dout[23] ) );
  DFFPOSX1 \myram/m14/d/d24/q_reg  ( .D(\myram/m14/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m14/dout[24] ) );
  DFFPOSX1 \myram/m14/d/d25/q_reg  ( .D(\myram/m14/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m14/dout[25] ) );
  DFFPOSX1 \myram/m14/d/d26/q_reg  ( .D(\myram/m14/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m14/dout[26] ) );
  DFFPOSX1 \myram/m14/d/d27/q_reg  ( .D(\myram/m14/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m14/dout[27] ) );
  DFFPOSX1 \myram/m14/d/d28/q_reg  ( .D(\myram/m14/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m14/dout[28] ) );
  DFFPOSX1 \myram/m14/d/d29/q_reg  ( .D(\myram/m14/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m14/dout[29] ) );
  DFFPOSX1 \myram/m14/d/d30/q_reg  ( .D(\myram/m14/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m14/dout[30] ) );
  DFFPOSX1 \myram/m14/d/d31/q_reg  ( .D(\myram/m14/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m14/dout[31] ) );
  DFFPOSX1 \myram/m13/d/d0/q_reg  ( .D(\myram/m13/mux_out[0] ), .CLK(clk), .Q(
        \myram/m13/dout[0] ) );
  DFFPOSX1 \myram/m13/d/d1/q_reg  ( .D(\myram/m13/mux_out[1] ), .CLK(clk), .Q(
        \myram/m13/dout[1] ) );
  DFFPOSX1 \myram/m13/d/d2/q_reg  ( .D(\myram/m13/mux_out[2] ), .CLK(clk), .Q(
        \myram/m13/dout[2] ) );
  DFFPOSX1 \myram/m13/d/d3/q_reg  ( .D(\myram/m13/mux_out[3] ), .CLK(clk), .Q(
        \myram/m13/dout[3] ) );
  DFFPOSX1 \myram/m13/d/d4/q_reg  ( .D(\myram/m13/mux_out[4] ), .CLK(clk), .Q(
        \myram/m13/dout[4] ) );
  DFFPOSX1 \myram/m13/d/d5/q_reg  ( .D(\myram/m13/mux_out[5] ), .CLK(clk), .Q(
        \myram/m13/dout[5] ) );
  DFFPOSX1 \myram/m13/d/d6/q_reg  ( .D(\myram/m13/mux_out[6] ), .CLK(clk), .Q(
        \myram/m13/dout[6] ) );
  DFFPOSX1 \myram/m13/d/d7/q_reg  ( .D(\myram/m13/mux_out[7] ), .CLK(clk), .Q(
        \myram/m13/dout[7] ) );
  DFFPOSX1 \myram/m13/d/d8/q_reg  ( .D(\myram/m13/mux_out[8] ), .CLK(clk), .Q(
        \myram/m13/dout[8] ) );
  DFFPOSX1 \myram/m13/d/d9/q_reg  ( .D(\myram/m13/mux_out[9] ), .CLK(clk), .Q(
        \myram/m13/dout[9] ) );
  DFFPOSX1 \myram/m13/d/d10/q_reg  ( .D(\myram/m13/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m13/dout[10] ) );
  DFFPOSX1 \myram/m13/d/d11/q_reg  ( .D(\myram/m13/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m13/dout[11] ) );
  DFFPOSX1 \myram/m13/d/d12/q_reg  ( .D(\myram/m13/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m13/dout[12] ) );
  DFFPOSX1 \myram/m13/d/d13/q_reg  ( .D(\myram/m13/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m13/dout[13] ) );
  DFFPOSX1 \myram/m13/d/d14/q_reg  ( .D(\myram/m13/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m13/dout[14] ) );
  DFFPOSX1 \myram/m13/d/d15/q_reg  ( .D(\myram/m13/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m13/dout[15] ) );
  DFFPOSX1 \myram/m13/d/d16/q_reg  ( .D(\myram/m13/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m13/dout[16] ) );
  DFFPOSX1 \myram/m13/d/d17/q_reg  ( .D(\myram/m13/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m13/dout[17] ) );
  DFFPOSX1 \myram/m13/d/d18/q_reg  ( .D(\myram/m13/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m13/dout[18] ) );
  DFFPOSX1 \myram/m13/d/d19/q_reg  ( .D(\myram/m13/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m13/dout[19] ) );
  DFFPOSX1 \myram/m13/d/d20/q_reg  ( .D(\myram/m13/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m13/dout[20] ) );
  DFFPOSX1 \myram/m13/d/d21/q_reg  ( .D(\myram/m13/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m13/dout[21] ) );
  DFFPOSX1 \myram/m13/d/d22/q_reg  ( .D(\myram/m13/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m13/dout[22] ) );
  DFFPOSX1 \myram/m13/d/d23/q_reg  ( .D(\myram/m13/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m13/dout[23] ) );
  DFFPOSX1 \myram/m13/d/d24/q_reg  ( .D(\myram/m13/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m13/dout[24] ) );
  DFFPOSX1 \myram/m13/d/d25/q_reg  ( .D(\myram/m13/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m13/dout[25] ) );
  DFFPOSX1 \myram/m13/d/d26/q_reg  ( .D(\myram/m13/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m13/dout[26] ) );
  DFFPOSX1 \myram/m13/d/d27/q_reg  ( .D(\myram/m13/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m13/dout[27] ) );
  DFFPOSX1 \myram/m13/d/d28/q_reg  ( .D(\myram/m13/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m13/dout[28] ) );
  DFFPOSX1 \myram/m13/d/d29/q_reg  ( .D(\myram/m13/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m13/dout[29] ) );
  DFFPOSX1 \myram/m13/d/d30/q_reg  ( .D(\myram/m13/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m13/dout[30] ) );
  DFFPOSX1 \myram/m13/d/d31/q_reg  ( .D(\myram/m13/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m13/dout[31] ) );
  DFFPOSX1 \myram/m12/d/d0/q_reg  ( .D(\myram/m12/mux_out[0] ), .CLK(clk), .Q(
        \myram/m12/dout[0] ) );
  DFFPOSX1 \myram/m12/d/d1/q_reg  ( .D(\myram/m12/mux_out[1] ), .CLK(clk), .Q(
        \myram/m12/dout[1] ) );
  DFFPOSX1 \myram/m12/d/d2/q_reg  ( .D(\myram/m12/mux_out[2] ), .CLK(clk), .Q(
        \myram/m12/dout[2] ) );
  DFFPOSX1 \myram/m12/d/d3/q_reg  ( .D(\myram/m12/mux_out[3] ), .CLK(clk), .Q(
        \myram/m12/dout[3] ) );
  DFFPOSX1 \myram/m12/d/d4/q_reg  ( .D(\myram/m12/mux_out[4] ), .CLK(clk), .Q(
        \myram/m12/dout[4] ) );
  DFFPOSX1 \myram/m12/d/d5/q_reg  ( .D(\myram/m12/mux_out[5] ), .CLK(clk), .Q(
        \myram/m12/dout[5] ) );
  DFFPOSX1 \myram/m12/d/d6/q_reg  ( .D(\myram/m12/mux_out[6] ), .CLK(clk), .Q(
        \myram/m12/dout[6] ) );
  DFFPOSX1 \myram/m12/d/d7/q_reg  ( .D(\myram/m12/mux_out[7] ), .CLK(clk), .Q(
        \myram/m12/dout[7] ) );
  DFFPOSX1 \myram/m12/d/d8/q_reg  ( .D(\myram/m12/mux_out[8] ), .CLK(clk), .Q(
        \myram/m12/dout[8] ) );
  DFFPOSX1 \myram/m12/d/d9/q_reg  ( .D(\myram/m12/mux_out[9] ), .CLK(clk), .Q(
        \myram/m12/dout[9] ) );
  DFFPOSX1 \myram/m12/d/d10/q_reg  ( .D(\myram/m12/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m12/dout[10] ) );
  DFFPOSX1 \myram/m12/d/d11/q_reg  ( .D(\myram/m12/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m12/dout[11] ) );
  DFFPOSX1 \myram/m12/d/d12/q_reg  ( .D(\myram/m12/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m12/dout[12] ) );
  DFFPOSX1 \myram/m12/d/d13/q_reg  ( .D(\myram/m12/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m12/dout[13] ) );
  DFFPOSX1 \myram/m12/d/d14/q_reg  ( .D(\myram/m12/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m12/dout[14] ) );
  DFFPOSX1 \myram/m12/d/d15/q_reg  ( .D(\myram/m12/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m12/dout[15] ) );
  DFFPOSX1 \myram/m12/d/d16/q_reg  ( .D(\myram/m12/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m12/dout[16] ) );
  DFFPOSX1 \myram/m12/d/d17/q_reg  ( .D(\myram/m12/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m12/dout[17] ) );
  DFFPOSX1 \myram/m12/d/d18/q_reg  ( .D(\myram/m12/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m12/dout[18] ) );
  DFFPOSX1 \myram/m12/d/d19/q_reg  ( .D(\myram/m12/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m12/dout[19] ) );
  DFFPOSX1 \myram/m12/d/d20/q_reg  ( .D(\myram/m12/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m12/dout[20] ) );
  DFFPOSX1 \myram/m12/d/d21/q_reg  ( .D(\myram/m12/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m12/dout[21] ) );
  DFFPOSX1 \myram/m12/d/d22/q_reg  ( .D(\myram/m12/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m12/dout[22] ) );
  DFFPOSX1 \myram/m12/d/d23/q_reg  ( .D(\myram/m12/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m12/dout[23] ) );
  DFFPOSX1 \myram/m12/d/d24/q_reg  ( .D(\myram/m12/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m12/dout[24] ) );
  DFFPOSX1 \myram/m12/d/d25/q_reg  ( .D(\myram/m12/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m12/dout[25] ) );
  DFFPOSX1 \myram/m12/d/d26/q_reg  ( .D(\myram/m12/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m12/dout[26] ) );
  DFFPOSX1 \myram/m12/d/d27/q_reg  ( .D(\myram/m12/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m12/dout[27] ) );
  DFFPOSX1 \myram/m12/d/d28/q_reg  ( .D(\myram/m12/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m12/dout[28] ) );
  DFFPOSX1 \myram/m12/d/d29/q_reg  ( .D(\myram/m12/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m12/dout[29] ) );
  DFFPOSX1 \myram/m12/d/d30/q_reg  ( .D(\myram/m12/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m12/dout[30] ) );
  DFFPOSX1 \myram/m12/d/d31/q_reg  ( .D(\myram/m12/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m12/dout[31] ) );
  DFFPOSX1 \myram/m11/d/d0/q_reg  ( .D(\myram/m11/mux_out[0] ), .CLK(clk), .Q(
        \myram/m11/dout[0] ) );
  DFFPOSX1 \myram/m11/d/d1/q_reg  ( .D(\myram/m11/mux_out[1] ), .CLK(clk), .Q(
        \myram/m11/dout[1] ) );
  DFFPOSX1 \myram/m11/d/d2/q_reg  ( .D(\myram/m11/mux_out[2] ), .CLK(clk), .Q(
        \myram/m11/dout[2] ) );
  DFFPOSX1 \myram/m11/d/d3/q_reg  ( .D(\myram/m11/mux_out[3] ), .CLK(clk), .Q(
        \myram/m11/dout[3] ) );
  DFFPOSX1 \myram/m11/d/d4/q_reg  ( .D(\myram/m11/mux_out[4] ), .CLK(clk), .Q(
        \myram/m11/dout[4] ) );
  DFFPOSX1 \myram/m11/d/d5/q_reg  ( .D(\myram/m11/mux_out[5] ), .CLK(clk), .Q(
        \myram/m11/dout[5] ) );
  DFFPOSX1 \myram/m11/d/d6/q_reg  ( .D(\myram/m11/mux_out[6] ), .CLK(clk), .Q(
        \myram/m11/dout[6] ) );
  DFFPOSX1 \myram/m11/d/d7/q_reg  ( .D(\myram/m11/mux_out[7] ), .CLK(clk), .Q(
        \myram/m11/dout[7] ) );
  DFFPOSX1 \myram/m11/d/d8/q_reg  ( .D(\myram/m11/mux_out[8] ), .CLK(clk), .Q(
        \myram/m11/dout[8] ) );
  DFFPOSX1 \myram/m11/d/d9/q_reg  ( .D(\myram/m11/mux_out[9] ), .CLK(clk), .Q(
        \myram/m11/dout[9] ) );
  DFFPOSX1 \myram/m11/d/d10/q_reg  ( .D(\myram/m11/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m11/dout[10] ) );
  DFFPOSX1 \myram/m11/d/d11/q_reg  ( .D(\myram/m11/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m11/dout[11] ) );
  DFFPOSX1 \myram/m11/d/d12/q_reg  ( .D(\myram/m11/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m11/dout[12] ) );
  DFFPOSX1 \myram/m11/d/d13/q_reg  ( .D(\myram/m11/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m11/dout[13] ) );
  DFFPOSX1 \myram/m11/d/d14/q_reg  ( .D(\myram/m11/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m11/dout[14] ) );
  DFFPOSX1 \myram/m11/d/d15/q_reg  ( .D(\myram/m11/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m11/dout[15] ) );
  DFFPOSX1 \myram/m11/d/d16/q_reg  ( .D(\myram/m11/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m11/dout[16] ) );
  DFFPOSX1 \myram/m11/d/d17/q_reg  ( .D(\myram/m11/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m11/dout[17] ) );
  DFFPOSX1 \myram/m11/d/d18/q_reg  ( .D(\myram/m11/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m11/dout[18] ) );
  DFFPOSX1 \myram/m11/d/d19/q_reg  ( .D(\myram/m11/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m11/dout[19] ) );
  DFFPOSX1 \myram/m11/d/d20/q_reg  ( .D(\myram/m11/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m11/dout[20] ) );
  DFFPOSX1 \myram/m11/d/d21/q_reg  ( .D(\myram/m11/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m11/dout[21] ) );
  DFFPOSX1 \myram/m11/d/d22/q_reg  ( .D(\myram/m11/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m11/dout[22] ) );
  DFFPOSX1 \myram/m11/d/d23/q_reg  ( .D(\myram/m11/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m11/dout[23] ) );
  DFFPOSX1 \myram/m11/d/d24/q_reg  ( .D(\myram/m11/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m11/dout[24] ) );
  DFFPOSX1 \myram/m11/d/d25/q_reg  ( .D(\myram/m11/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m11/dout[25] ) );
  DFFPOSX1 \myram/m11/d/d26/q_reg  ( .D(\myram/m11/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m11/dout[26] ) );
  DFFPOSX1 \myram/m11/d/d27/q_reg  ( .D(\myram/m11/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m11/dout[27] ) );
  DFFPOSX1 \myram/m11/d/d28/q_reg  ( .D(\myram/m11/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m11/dout[28] ) );
  DFFPOSX1 \myram/m11/d/d29/q_reg  ( .D(\myram/m11/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m11/dout[29] ) );
  DFFPOSX1 \myram/m11/d/d30/q_reg  ( .D(\myram/m11/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m11/dout[30] ) );
  DFFPOSX1 \myram/m11/d/d31/q_reg  ( .D(\myram/m11/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m11/dout[31] ) );
  DFFPOSX1 \myram/m10/d/d0/q_reg  ( .D(\myram/m10/mux_out[0] ), .CLK(clk), .Q(
        \myram/m10/dout[0] ) );
  DFFPOSX1 \myram/m10/d/d1/q_reg  ( .D(\myram/m10/mux_out[1] ), .CLK(clk), .Q(
        \myram/m10/dout[1] ) );
  DFFPOSX1 \myram/m10/d/d2/q_reg  ( .D(\myram/m10/mux_out[2] ), .CLK(clk), .Q(
        \myram/m10/dout[2] ) );
  DFFPOSX1 \myram/m10/d/d3/q_reg  ( .D(\myram/m10/mux_out[3] ), .CLK(clk), .Q(
        \myram/m10/dout[3] ) );
  DFFPOSX1 \myram/m10/d/d4/q_reg  ( .D(\myram/m10/mux_out[4] ), .CLK(clk), .Q(
        \myram/m10/dout[4] ) );
  DFFPOSX1 \myram/m10/d/d5/q_reg  ( .D(\myram/m10/mux_out[5] ), .CLK(clk), .Q(
        \myram/m10/dout[5] ) );
  DFFPOSX1 \myram/m10/d/d6/q_reg  ( .D(\myram/m10/mux_out[6] ), .CLK(clk), .Q(
        \myram/m10/dout[6] ) );
  DFFPOSX1 \myram/m10/d/d7/q_reg  ( .D(\myram/m10/mux_out[7] ), .CLK(clk), .Q(
        \myram/m10/dout[7] ) );
  DFFPOSX1 \myram/m10/d/d8/q_reg  ( .D(\myram/m10/mux_out[8] ), .CLK(clk), .Q(
        \myram/m10/dout[8] ) );
  DFFPOSX1 \myram/m10/d/d9/q_reg  ( .D(\myram/m10/mux_out[9] ), .CLK(clk), .Q(
        \myram/m10/dout[9] ) );
  DFFPOSX1 \myram/m10/d/d10/q_reg  ( .D(\myram/m10/mux_out[10] ), .CLK(clk), 
        .Q(\myram/m10/dout[10] ) );
  DFFPOSX1 \myram/m10/d/d11/q_reg  ( .D(\myram/m10/mux_out[11] ), .CLK(clk), 
        .Q(\myram/m10/dout[11] ) );
  DFFPOSX1 \myram/m10/d/d12/q_reg  ( .D(\myram/m10/mux_out[12] ), .CLK(clk), 
        .Q(\myram/m10/dout[12] ) );
  DFFPOSX1 \myram/m10/d/d13/q_reg  ( .D(\myram/m10/mux_out[13] ), .CLK(clk), 
        .Q(\myram/m10/dout[13] ) );
  DFFPOSX1 \myram/m10/d/d14/q_reg  ( .D(\myram/m10/mux_out[14] ), .CLK(clk), 
        .Q(\myram/m10/dout[14] ) );
  DFFPOSX1 \myram/m10/d/d15/q_reg  ( .D(\myram/m10/mux_out[15] ), .CLK(clk), 
        .Q(\myram/m10/dout[15] ) );
  DFFPOSX1 \myram/m10/d/d16/q_reg  ( .D(\myram/m10/mux_out[16] ), .CLK(clk), 
        .Q(\myram/m10/dout[16] ) );
  DFFPOSX1 \myram/m10/d/d17/q_reg  ( .D(\myram/m10/mux_out[17] ), .CLK(clk), 
        .Q(\myram/m10/dout[17] ) );
  DFFPOSX1 \myram/m10/d/d18/q_reg  ( .D(\myram/m10/mux_out[18] ), .CLK(clk), 
        .Q(\myram/m10/dout[18] ) );
  DFFPOSX1 \myram/m10/d/d19/q_reg  ( .D(\myram/m10/mux_out[19] ), .CLK(clk), 
        .Q(\myram/m10/dout[19] ) );
  DFFPOSX1 \myram/m10/d/d20/q_reg  ( .D(\myram/m10/mux_out[20] ), .CLK(clk), 
        .Q(\myram/m10/dout[20] ) );
  DFFPOSX1 \myram/m10/d/d21/q_reg  ( .D(\myram/m10/mux_out[21] ), .CLK(clk), 
        .Q(\myram/m10/dout[21] ) );
  DFFPOSX1 \myram/m10/d/d22/q_reg  ( .D(\myram/m10/mux_out[22] ), .CLK(clk), 
        .Q(\myram/m10/dout[22] ) );
  DFFPOSX1 \myram/m10/d/d23/q_reg  ( .D(\myram/m10/mux_out[23] ), .CLK(clk), 
        .Q(\myram/m10/dout[23] ) );
  DFFPOSX1 \myram/m10/d/d24/q_reg  ( .D(\myram/m10/mux_out[24] ), .CLK(clk), 
        .Q(\myram/m10/dout[24] ) );
  DFFPOSX1 \myram/m10/d/d25/q_reg  ( .D(\myram/m10/mux_out[25] ), .CLK(clk), 
        .Q(\myram/m10/dout[25] ) );
  DFFPOSX1 \myram/m10/d/d26/q_reg  ( .D(\myram/m10/mux_out[26] ), .CLK(clk), 
        .Q(\myram/m10/dout[26] ) );
  DFFPOSX1 \myram/m10/d/d27/q_reg  ( .D(\myram/m10/mux_out[27] ), .CLK(clk), 
        .Q(\myram/m10/dout[27] ) );
  DFFPOSX1 \myram/m10/d/d28/q_reg  ( .D(\myram/m10/mux_out[28] ), .CLK(clk), 
        .Q(\myram/m10/dout[28] ) );
  DFFPOSX1 \myram/m10/d/d29/q_reg  ( .D(\myram/m10/mux_out[29] ), .CLK(clk), 
        .Q(\myram/m10/dout[29] ) );
  DFFPOSX1 \myram/m10/d/d30/q_reg  ( .D(\myram/m10/mux_out[30] ), .CLK(clk), 
        .Q(\myram/m10/dout[30] ) );
  DFFPOSX1 \myram/m10/d/d31/q_reg  ( .D(\myram/m10/mux_out[31] ), .CLK(clk), 
        .Q(\myram/m10/dout[31] ) );
  DFFPOSX1 \myram/m9/d/d0/q_reg  ( .D(\myram/m9/mux_out[0] ), .CLK(clk), .Q(
        \myram/m9/dout[0] ) );
  DFFPOSX1 \myram/m9/d/d1/q_reg  ( .D(\myram/m9/mux_out[1] ), .CLK(clk), .Q(
        \myram/m9/dout[1] ) );
  DFFPOSX1 \myram/m9/d/d2/q_reg  ( .D(\myram/m9/mux_out[2] ), .CLK(clk), .Q(
        \myram/m9/dout[2] ) );
  DFFPOSX1 \myram/m9/d/d3/q_reg  ( .D(\myram/m9/mux_out[3] ), .CLK(clk), .Q(
        \myram/m9/dout[3] ) );
  DFFPOSX1 \myram/m9/d/d4/q_reg  ( .D(\myram/m9/mux_out[4] ), .CLK(clk), .Q(
        \myram/m9/dout[4] ) );
  DFFPOSX1 \myram/m9/d/d5/q_reg  ( .D(\myram/m9/mux_out[5] ), .CLK(clk), .Q(
        \myram/m9/dout[5] ) );
  DFFPOSX1 \myram/m9/d/d6/q_reg  ( .D(\myram/m9/mux_out[6] ), .CLK(clk), .Q(
        \myram/m9/dout[6] ) );
  DFFPOSX1 \myram/m9/d/d7/q_reg  ( .D(\myram/m9/mux_out[7] ), .CLK(clk), .Q(
        \myram/m9/dout[7] ) );
  DFFPOSX1 \myram/m9/d/d8/q_reg  ( .D(\myram/m9/mux_out[8] ), .CLK(clk), .Q(
        \myram/m9/dout[8] ) );
  DFFPOSX1 \myram/m9/d/d9/q_reg  ( .D(\myram/m9/mux_out[9] ), .CLK(clk), .Q(
        \myram/m9/dout[9] ) );
  DFFPOSX1 \myram/m9/d/d10/q_reg  ( .D(\myram/m9/mux_out[10] ), .CLK(clk), .Q(
        \myram/m9/dout[10] ) );
  DFFPOSX1 \myram/m9/d/d11/q_reg  ( .D(\myram/m9/mux_out[11] ), .CLK(clk), .Q(
        \myram/m9/dout[11] ) );
  DFFPOSX1 \myram/m9/d/d12/q_reg  ( .D(\myram/m9/mux_out[12] ), .CLK(clk), .Q(
        \myram/m9/dout[12] ) );
  DFFPOSX1 \myram/m9/d/d13/q_reg  ( .D(\myram/m9/mux_out[13] ), .CLK(clk), .Q(
        \myram/m9/dout[13] ) );
  DFFPOSX1 \myram/m9/d/d14/q_reg  ( .D(\myram/m9/mux_out[14] ), .CLK(clk), .Q(
        \myram/m9/dout[14] ) );
  DFFPOSX1 \myram/m9/d/d15/q_reg  ( .D(\myram/m9/mux_out[15] ), .CLK(clk), .Q(
        \myram/m9/dout[15] ) );
  DFFPOSX1 \myram/m9/d/d16/q_reg  ( .D(\myram/m9/mux_out[16] ), .CLK(clk), .Q(
        \myram/m9/dout[16] ) );
  DFFPOSX1 \myram/m9/d/d17/q_reg  ( .D(\myram/m9/mux_out[17] ), .CLK(clk), .Q(
        \myram/m9/dout[17] ) );
  DFFPOSX1 \myram/m9/d/d18/q_reg  ( .D(\myram/m9/mux_out[18] ), .CLK(clk), .Q(
        \myram/m9/dout[18] ) );
  DFFPOSX1 \myram/m9/d/d19/q_reg  ( .D(\myram/m9/mux_out[19] ), .CLK(clk), .Q(
        \myram/m9/dout[19] ) );
  DFFPOSX1 \myram/m9/d/d20/q_reg  ( .D(\myram/m9/mux_out[20] ), .CLK(clk), .Q(
        \myram/m9/dout[20] ) );
  DFFPOSX1 \myram/m9/d/d21/q_reg  ( .D(\myram/m9/mux_out[21] ), .CLK(clk), .Q(
        \myram/m9/dout[21] ) );
  DFFPOSX1 \myram/m9/d/d22/q_reg  ( .D(\myram/m9/mux_out[22] ), .CLK(clk), .Q(
        \myram/m9/dout[22] ) );
  DFFPOSX1 \myram/m9/d/d23/q_reg  ( .D(\myram/m9/mux_out[23] ), .CLK(clk), .Q(
        \myram/m9/dout[23] ) );
  DFFPOSX1 \myram/m9/d/d24/q_reg  ( .D(\myram/m9/mux_out[24] ), .CLK(clk), .Q(
        \myram/m9/dout[24] ) );
  DFFPOSX1 \myram/m9/d/d25/q_reg  ( .D(\myram/m9/mux_out[25] ), .CLK(clk), .Q(
        \myram/m9/dout[25] ) );
  DFFPOSX1 \myram/m9/d/d26/q_reg  ( .D(\myram/m9/mux_out[26] ), .CLK(clk), .Q(
        \myram/m9/dout[26] ) );
  DFFPOSX1 \myram/m9/d/d27/q_reg  ( .D(\myram/m9/mux_out[27] ), .CLK(clk), .Q(
        \myram/m9/dout[27] ) );
  DFFPOSX1 \myram/m9/d/d28/q_reg  ( .D(\myram/m9/mux_out[28] ), .CLK(clk), .Q(
        \myram/m9/dout[28] ) );
  DFFPOSX1 \myram/m9/d/d29/q_reg  ( .D(\myram/m9/mux_out[29] ), .CLK(clk), .Q(
        \myram/m9/dout[29] ) );
  DFFPOSX1 \myram/m9/d/d30/q_reg  ( .D(\myram/m9/mux_out[30] ), .CLK(clk), .Q(
        \myram/m9/dout[30] ) );
  DFFPOSX1 \myram/m9/d/d31/q_reg  ( .D(\myram/m9/mux_out[31] ), .CLK(clk), .Q(
        \myram/m9/dout[31] ) );
  DFFPOSX1 \myram/m8/d/d0/q_reg  ( .D(\myram/m8/mux_out[0] ), .CLK(clk), .Q(
        \myram/m8/dout[0] ) );
  DFFPOSX1 \myram/m8/d/d1/q_reg  ( .D(\myram/m8/mux_out[1] ), .CLK(clk), .Q(
        \myram/m8/dout[1] ) );
  DFFPOSX1 \myram/m8/d/d2/q_reg  ( .D(\myram/m8/mux_out[2] ), .CLK(clk), .Q(
        \myram/m8/dout[2] ) );
  DFFPOSX1 \myram/m8/d/d3/q_reg  ( .D(\myram/m8/mux_out[3] ), .CLK(clk), .Q(
        \myram/m8/dout[3] ) );
  DFFPOSX1 \myram/m8/d/d4/q_reg  ( .D(\myram/m8/mux_out[4] ), .CLK(clk), .Q(
        \myram/m8/dout[4] ) );
  DFFPOSX1 \myram/m8/d/d5/q_reg  ( .D(\myram/m8/mux_out[5] ), .CLK(clk), .Q(
        \myram/m8/dout[5] ) );
  DFFPOSX1 \myram/m8/d/d6/q_reg  ( .D(\myram/m8/mux_out[6] ), .CLK(clk), .Q(
        \myram/m8/dout[6] ) );
  DFFPOSX1 \myram/m8/d/d7/q_reg  ( .D(\myram/m8/mux_out[7] ), .CLK(clk), .Q(
        \myram/m8/dout[7] ) );
  DFFPOSX1 \myram/m8/d/d8/q_reg  ( .D(\myram/m8/mux_out[8] ), .CLK(clk), .Q(
        \myram/m8/dout[8] ) );
  DFFPOSX1 \myram/m8/d/d9/q_reg  ( .D(\myram/m8/mux_out[9] ), .CLK(clk), .Q(
        \myram/m8/dout[9] ) );
  DFFPOSX1 \myram/m8/d/d10/q_reg  ( .D(\myram/m8/mux_out[10] ), .CLK(clk), .Q(
        \myram/m8/dout[10] ) );
  DFFPOSX1 \myram/m8/d/d11/q_reg  ( .D(\myram/m8/mux_out[11] ), .CLK(clk), .Q(
        \myram/m8/dout[11] ) );
  DFFPOSX1 \myram/m8/d/d12/q_reg  ( .D(\myram/m8/mux_out[12] ), .CLK(clk), .Q(
        \myram/m8/dout[12] ) );
  DFFPOSX1 \myram/m8/d/d13/q_reg  ( .D(\myram/m8/mux_out[13] ), .CLK(clk), .Q(
        \myram/m8/dout[13] ) );
  DFFPOSX1 \myram/m8/d/d14/q_reg  ( .D(\myram/m8/mux_out[14] ), .CLK(clk), .Q(
        \myram/m8/dout[14] ) );
  DFFPOSX1 \myram/m8/d/d15/q_reg  ( .D(\myram/m8/mux_out[15] ), .CLK(clk), .Q(
        \myram/m8/dout[15] ) );
  DFFPOSX1 \myram/m8/d/d16/q_reg  ( .D(\myram/m8/mux_out[16] ), .CLK(clk), .Q(
        \myram/m8/dout[16] ) );
  DFFPOSX1 \myram/m8/d/d17/q_reg  ( .D(\myram/m8/mux_out[17] ), .CLK(clk), .Q(
        \myram/m8/dout[17] ) );
  DFFPOSX1 \myram/m8/d/d18/q_reg  ( .D(\myram/m8/mux_out[18] ), .CLK(clk), .Q(
        \myram/m8/dout[18] ) );
  DFFPOSX1 \myram/m8/d/d19/q_reg  ( .D(\myram/m8/mux_out[19] ), .CLK(clk), .Q(
        \myram/m8/dout[19] ) );
  DFFPOSX1 \myram/m8/d/d20/q_reg  ( .D(\myram/m8/mux_out[20] ), .CLK(clk), .Q(
        \myram/m8/dout[20] ) );
  DFFPOSX1 \myram/m8/d/d21/q_reg  ( .D(\myram/m8/mux_out[21] ), .CLK(clk), .Q(
        \myram/m8/dout[21] ) );
  DFFPOSX1 \myram/m8/d/d22/q_reg  ( .D(\myram/m8/mux_out[22] ), .CLK(clk), .Q(
        \myram/m8/dout[22] ) );
  DFFPOSX1 \myram/m8/d/d23/q_reg  ( .D(\myram/m8/mux_out[23] ), .CLK(clk), .Q(
        \myram/m8/dout[23] ) );
  DFFPOSX1 \myram/m8/d/d24/q_reg  ( .D(\myram/m8/mux_out[24] ), .CLK(clk), .Q(
        \myram/m8/dout[24] ) );
  DFFPOSX1 \myram/m8/d/d25/q_reg  ( .D(\myram/m8/mux_out[25] ), .CLK(clk), .Q(
        \myram/m8/dout[25] ) );
  DFFPOSX1 \myram/m8/d/d26/q_reg  ( .D(\myram/m8/mux_out[26] ), .CLK(clk), .Q(
        \myram/m8/dout[26] ) );
  DFFPOSX1 \myram/m8/d/d27/q_reg  ( .D(\myram/m8/mux_out[27] ), .CLK(clk), .Q(
        \myram/m8/dout[27] ) );
  DFFPOSX1 \myram/m8/d/d28/q_reg  ( .D(\myram/m8/mux_out[28] ), .CLK(clk), .Q(
        \myram/m8/dout[28] ) );
  DFFPOSX1 \myram/m8/d/d29/q_reg  ( .D(\myram/m8/mux_out[29] ), .CLK(clk), .Q(
        \myram/m8/dout[29] ) );
  DFFPOSX1 \myram/m8/d/d30/q_reg  ( .D(\myram/m8/mux_out[30] ), .CLK(clk), .Q(
        \myram/m8/dout[30] ) );
  DFFPOSX1 \myram/m8/d/d31/q_reg  ( .D(\myram/m8/mux_out[31] ), .CLK(clk), .Q(
        \myram/m8/dout[31] ) );
  DFFPOSX1 \myram/m7/d/d0/q_reg  ( .D(\myram/m7/mux_out[0] ), .CLK(clk), .Q(
        \myram/m7/dout[0] ) );
  DFFPOSX1 \myram/m7/d/d1/q_reg  ( .D(\myram/m7/mux_out[1] ), .CLK(clk), .Q(
        \myram/m7/dout[1] ) );
  DFFPOSX1 \myram/m7/d/d2/q_reg  ( .D(\myram/m7/mux_out[2] ), .CLK(clk), .Q(
        \myram/m7/dout[2] ) );
  DFFPOSX1 \myram/m7/d/d3/q_reg  ( .D(\myram/m7/mux_out[3] ), .CLK(clk), .Q(
        \myram/m7/dout[3] ) );
  DFFPOSX1 \myram/m7/d/d4/q_reg  ( .D(\myram/m7/mux_out[4] ), .CLK(clk), .Q(
        \myram/m7/dout[4] ) );
  DFFPOSX1 \myram/m7/d/d5/q_reg  ( .D(\myram/m7/mux_out[5] ), .CLK(clk), .Q(
        \myram/m7/dout[5] ) );
  DFFPOSX1 \myram/m7/d/d6/q_reg  ( .D(\myram/m7/mux_out[6] ), .CLK(clk), .Q(
        \myram/m7/dout[6] ) );
  DFFPOSX1 \myram/m7/d/d7/q_reg  ( .D(\myram/m7/mux_out[7] ), .CLK(clk), .Q(
        \myram/m7/dout[7] ) );
  DFFPOSX1 \myram/m7/d/d8/q_reg  ( .D(\myram/m7/mux_out[8] ), .CLK(clk), .Q(
        \myram/m7/dout[8] ) );
  DFFPOSX1 \myram/m7/d/d9/q_reg  ( .D(\myram/m7/mux_out[9] ), .CLK(clk), .Q(
        \myram/m7/dout[9] ) );
  DFFPOSX1 \myram/m7/d/d10/q_reg  ( .D(\myram/m7/mux_out[10] ), .CLK(clk), .Q(
        \myram/m7/dout[10] ) );
  DFFPOSX1 \myram/m7/d/d11/q_reg  ( .D(\myram/m7/mux_out[11] ), .CLK(clk), .Q(
        \myram/m7/dout[11] ) );
  DFFPOSX1 \myram/m7/d/d12/q_reg  ( .D(\myram/m7/mux_out[12] ), .CLK(clk), .Q(
        \myram/m7/dout[12] ) );
  DFFPOSX1 \myram/m7/d/d13/q_reg  ( .D(\myram/m7/mux_out[13] ), .CLK(clk), .Q(
        \myram/m7/dout[13] ) );
  DFFPOSX1 \myram/m7/d/d14/q_reg  ( .D(\myram/m7/mux_out[14] ), .CLK(clk), .Q(
        \myram/m7/dout[14] ) );
  DFFPOSX1 \myram/m7/d/d15/q_reg  ( .D(\myram/m7/mux_out[15] ), .CLK(clk), .Q(
        \myram/m7/dout[15] ) );
  DFFPOSX1 \myram/m7/d/d16/q_reg  ( .D(\myram/m7/mux_out[16] ), .CLK(clk), .Q(
        \myram/m7/dout[16] ) );
  DFFPOSX1 \myram/m7/d/d17/q_reg  ( .D(\myram/m7/mux_out[17] ), .CLK(clk), .Q(
        \myram/m7/dout[17] ) );
  DFFPOSX1 \myram/m7/d/d18/q_reg  ( .D(\myram/m7/mux_out[18] ), .CLK(clk), .Q(
        \myram/m7/dout[18] ) );
  DFFPOSX1 \myram/m7/d/d19/q_reg  ( .D(\myram/m7/mux_out[19] ), .CLK(clk), .Q(
        \myram/m7/dout[19] ) );
  DFFPOSX1 \myram/m7/d/d20/q_reg  ( .D(\myram/m7/mux_out[20] ), .CLK(clk), .Q(
        \myram/m7/dout[20] ) );
  DFFPOSX1 \myram/m7/d/d21/q_reg  ( .D(\myram/m7/mux_out[21] ), .CLK(clk), .Q(
        \myram/m7/dout[21] ) );
  DFFPOSX1 \myram/m7/d/d22/q_reg  ( .D(\myram/m7/mux_out[22] ), .CLK(clk), .Q(
        \myram/m7/dout[22] ) );
  DFFPOSX1 \myram/m7/d/d23/q_reg  ( .D(\myram/m7/mux_out[23] ), .CLK(clk), .Q(
        \myram/m7/dout[23] ) );
  DFFPOSX1 \myram/m7/d/d24/q_reg  ( .D(\myram/m7/mux_out[24] ), .CLK(clk), .Q(
        \myram/m7/dout[24] ) );
  DFFPOSX1 \myram/m7/d/d25/q_reg  ( .D(\myram/m7/mux_out[25] ), .CLK(clk), .Q(
        \myram/m7/dout[25] ) );
  DFFPOSX1 \myram/m7/d/d26/q_reg  ( .D(\myram/m7/mux_out[26] ), .CLK(clk), .Q(
        \myram/m7/dout[26] ) );
  DFFPOSX1 \myram/m7/d/d27/q_reg  ( .D(\myram/m7/mux_out[27] ), .CLK(clk), .Q(
        \myram/m7/dout[27] ) );
  DFFPOSX1 \myram/m7/d/d28/q_reg  ( .D(\myram/m7/mux_out[28] ), .CLK(clk), .Q(
        \myram/m7/dout[28] ) );
  DFFPOSX1 \myram/m7/d/d29/q_reg  ( .D(\myram/m7/mux_out[29] ), .CLK(clk), .Q(
        \myram/m7/dout[29] ) );
  DFFPOSX1 \myram/m7/d/d30/q_reg  ( .D(\myram/m7/mux_out[30] ), .CLK(clk), .Q(
        \myram/m7/dout[30] ) );
  DFFPOSX1 \myram/m7/d/d31/q_reg  ( .D(\myram/m7/mux_out[31] ), .CLK(clk), .Q(
        \myram/m7/dout[31] ) );
  DFFPOSX1 \myram/m6/d/d0/q_reg  ( .D(\myram/m6/mux_out[0] ), .CLK(clk), .Q(
        \myram/m6/dout[0] ) );
  DFFPOSX1 \myram/m6/d/d1/q_reg  ( .D(\myram/m6/mux_out[1] ), .CLK(clk), .Q(
        \myram/m6/dout[1] ) );
  DFFPOSX1 \myram/m6/d/d2/q_reg  ( .D(\myram/m6/mux_out[2] ), .CLK(clk), .Q(
        \myram/m6/dout[2] ) );
  DFFPOSX1 \myram/m6/d/d3/q_reg  ( .D(\myram/m6/mux_out[3] ), .CLK(clk), .Q(
        \myram/m6/dout[3] ) );
  DFFPOSX1 \myram/m6/d/d4/q_reg  ( .D(\myram/m6/mux_out[4] ), .CLK(clk), .Q(
        \myram/m6/dout[4] ) );
  DFFPOSX1 \myram/m6/d/d5/q_reg  ( .D(\myram/m6/mux_out[5] ), .CLK(clk), .Q(
        \myram/m6/dout[5] ) );
  DFFPOSX1 \myram/m6/d/d6/q_reg  ( .D(\myram/m6/mux_out[6] ), .CLK(clk), .Q(
        \myram/m6/dout[6] ) );
  DFFPOSX1 \myram/m6/d/d7/q_reg  ( .D(\myram/m6/mux_out[7] ), .CLK(clk), .Q(
        \myram/m6/dout[7] ) );
  DFFPOSX1 \myram/m6/d/d8/q_reg  ( .D(\myram/m6/mux_out[8] ), .CLK(clk), .Q(
        \myram/m6/dout[8] ) );
  DFFPOSX1 \myram/m6/d/d9/q_reg  ( .D(\myram/m6/mux_out[9] ), .CLK(clk), .Q(
        \myram/m6/dout[9] ) );
  DFFPOSX1 \myram/m6/d/d10/q_reg  ( .D(\myram/m6/mux_out[10] ), .CLK(clk), .Q(
        \myram/m6/dout[10] ) );
  DFFPOSX1 \myram/m6/d/d11/q_reg  ( .D(\myram/m6/mux_out[11] ), .CLK(clk), .Q(
        \myram/m6/dout[11] ) );
  DFFPOSX1 \myram/m6/d/d12/q_reg  ( .D(\myram/m6/mux_out[12] ), .CLK(clk), .Q(
        \myram/m6/dout[12] ) );
  DFFPOSX1 \myram/m6/d/d13/q_reg  ( .D(\myram/m6/mux_out[13] ), .CLK(clk), .Q(
        \myram/m6/dout[13] ) );
  DFFPOSX1 \myram/m6/d/d14/q_reg  ( .D(\myram/m6/mux_out[14] ), .CLK(clk), .Q(
        \myram/m6/dout[14] ) );
  DFFPOSX1 \myram/m6/d/d15/q_reg  ( .D(\myram/m6/mux_out[15] ), .CLK(clk), .Q(
        \myram/m6/dout[15] ) );
  DFFPOSX1 \myram/m6/d/d16/q_reg  ( .D(\myram/m6/mux_out[16] ), .CLK(clk), .Q(
        \myram/m6/dout[16] ) );
  DFFPOSX1 \myram/m6/d/d17/q_reg  ( .D(\myram/m6/mux_out[17] ), .CLK(clk), .Q(
        \myram/m6/dout[17] ) );
  DFFPOSX1 \myram/m6/d/d18/q_reg  ( .D(\myram/m6/mux_out[18] ), .CLK(clk), .Q(
        \myram/m6/dout[18] ) );
  DFFPOSX1 \myram/m6/d/d19/q_reg  ( .D(\myram/m6/mux_out[19] ), .CLK(clk), .Q(
        \myram/m6/dout[19] ) );
  DFFPOSX1 \myram/m6/d/d20/q_reg  ( .D(\myram/m6/mux_out[20] ), .CLK(clk), .Q(
        \myram/m6/dout[20] ) );
  DFFPOSX1 \myram/m6/d/d21/q_reg  ( .D(\myram/m6/mux_out[21] ), .CLK(clk), .Q(
        \myram/m6/dout[21] ) );
  DFFPOSX1 \myram/m6/d/d22/q_reg  ( .D(\myram/m6/mux_out[22] ), .CLK(clk), .Q(
        \myram/m6/dout[22] ) );
  DFFPOSX1 \myram/m6/d/d23/q_reg  ( .D(\myram/m6/mux_out[23] ), .CLK(clk), .Q(
        \myram/m6/dout[23] ) );
  DFFPOSX1 \myram/m6/d/d24/q_reg  ( .D(\myram/m6/mux_out[24] ), .CLK(clk), .Q(
        \myram/m6/dout[24] ) );
  DFFPOSX1 \myram/m6/d/d25/q_reg  ( .D(\myram/m6/mux_out[25] ), .CLK(clk), .Q(
        \myram/m6/dout[25] ) );
  DFFPOSX1 \myram/m6/d/d26/q_reg  ( .D(\myram/m6/mux_out[26] ), .CLK(clk), .Q(
        \myram/m6/dout[26] ) );
  DFFPOSX1 \myram/m6/d/d27/q_reg  ( .D(\myram/m6/mux_out[27] ), .CLK(clk), .Q(
        \myram/m6/dout[27] ) );
  DFFPOSX1 \myram/m6/d/d28/q_reg  ( .D(\myram/m6/mux_out[28] ), .CLK(clk), .Q(
        \myram/m6/dout[28] ) );
  DFFPOSX1 \myram/m6/d/d29/q_reg  ( .D(\myram/m6/mux_out[29] ), .CLK(clk), .Q(
        \myram/m6/dout[29] ) );
  DFFPOSX1 \myram/m6/d/d30/q_reg  ( .D(\myram/m6/mux_out[30] ), .CLK(clk), .Q(
        \myram/m6/dout[30] ) );
  DFFPOSX1 \myram/m6/d/d31/q_reg  ( .D(\myram/m6/mux_out[31] ), .CLK(clk), .Q(
        \myram/m6/dout[31] ) );
  DFFPOSX1 \myram/m5/d/d0/q_reg  ( .D(\myram/m5/mux_out[0] ), .CLK(clk), .Q(
        \myram/m5/dout[0] ) );
  DFFPOSX1 \myram/m5/d/d1/q_reg  ( .D(\myram/m5/mux_out[1] ), .CLK(clk), .Q(
        \myram/m5/dout[1] ) );
  DFFPOSX1 \myram/m5/d/d2/q_reg  ( .D(\myram/m5/mux_out[2] ), .CLK(clk), .Q(
        \myram/m5/dout[2] ) );
  DFFPOSX1 \myram/m5/d/d3/q_reg  ( .D(\myram/m5/mux_out[3] ), .CLK(clk), .Q(
        \myram/m5/dout[3] ) );
  DFFPOSX1 \myram/m5/d/d4/q_reg  ( .D(\myram/m5/mux_out[4] ), .CLK(clk), .Q(
        \myram/m5/dout[4] ) );
  DFFPOSX1 \myram/m5/d/d5/q_reg  ( .D(\myram/m5/mux_out[5] ), .CLK(clk), .Q(
        \myram/m5/dout[5] ) );
  DFFPOSX1 \myram/m5/d/d6/q_reg  ( .D(\myram/m5/mux_out[6] ), .CLK(clk), .Q(
        \myram/m5/dout[6] ) );
  DFFPOSX1 \myram/m5/d/d7/q_reg  ( .D(\myram/m5/mux_out[7] ), .CLK(clk), .Q(
        \myram/m5/dout[7] ) );
  DFFPOSX1 \myram/m5/d/d8/q_reg  ( .D(\myram/m5/mux_out[8] ), .CLK(clk), .Q(
        \myram/m5/dout[8] ) );
  DFFPOSX1 \myram/m5/d/d9/q_reg  ( .D(\myram/m5/mux_out[9] ), .CLK(clk), .Q(
        \myram/m5/dout[9] ) );
  DFFPOSX1 \myram/m5/d/d10/q_reg  ( .D(\myram/m5/mux_out[10] ), .CLK(clk), .Q(
        \myram/m5/dout[10] ) );
  DFFPOSX1 \myram/m5/d/d11/q_reg  ( .D(\myram/m5/mux_out[11] ), .CLK(clk), .Q(
        \myram/m5/dout[11] ) );
  DFFPOSX1 \myram/m5/d/d12/q_reg  ( .D(\myram/m5/mux_out[12] ), .CLK(clk), .Q(
        \myram/m5/dout[12] ) );
  DFFPOSX1 \myram/m5/d/d13/q_reg  ( .D(\myram/m5/mux_out[13] ), .CLK(clk), .Q(
        \myram/m5/dout[13] ) );
  DFFPOSX1 \myram/m5/d/d14/q_reg  ( .D(\myram/m5/mux_out[14] ), .CLK(clk), .Q(
        \myram/m5/dout[14] ) );
  DFFPOSX1 \myram/m5/d/d15/q_reg  ( .D(\myram/m5/mux_out[15] ), .CLK(clk), .Q(
        \myram/m5/dout[15] ) );
  DFFPOSX1 \myram/m5/d/d16/q_reg  ( .D(\myram/m5/mux_out[16] ), .CLK(clk), .Q(
        \myram/m5/dout[16] ) );
  DFFPOSX1 \myram/m5/d/d17/q_reg  ( .D(\myram/m5/mux_out[17] ), .CLK(clk), .Q(
        \myram/m5/dout[17] ) );
  DFFPOSX1 \myram/m5/d/d18/q_reg  ( .D(\myram/m5/mux_out[18] ), .CLK(clk), .Q(
        \myram/m5/dout[18] ) );
  DFFPOSX1 \myram/m5/d/d19/q_reg  ( .D(\myram/m5/mux_out[19] ), .CLK(clk), .Q(
        \myram/m5/dout[19] ) );
  DFFPOSX1 \myram/m5/d/d20/q_reg  ( .D(\myram/m5/mux_out[20] ), .CLK(clk), .Q(
        \myram/m5/dout[20] ) );
  DFFPOSX1 \myram/m5/d/d21/q_reg  ( .D(\myram/m5/mux_out[21] ), .CLK(clk), .Q(
        \myram/m5/dout[21] ) );
  DFFPOSX1 \myram/m5/d/d22/q_reg  ( .D(\myram/m5/mux_out[22] ), .CLK(clk), .Q(
        \myram/m5/dout[22] ) );
  DFFPOSX1 \myram/m5/d/d23/q_reg  ( .D(\myram/m5/mux_out[23] ), .CLK(clk), .Q(
        \myram/m5/dout[23] ) );
  DFFPOSX1 \myram/m5/d/d24/q_reg  ( .D(\myram/m5/mux_out[24] ), .CLK(clk), .Q(
        \myram/m5/dout[24] ) );
  DFFPOSX1 \myram/m5/d/d25/q_reg  ( .D(\myram/m5/mux_out[25] ), .CLK(clk), .Q(
        \myram/m5/dout[25] ) );
  DFFPOSX1 \myram/m5/d/d26/q_reg  ( .D(\myram/m5/mux_out[26] ), .CLK(clk), .Q(
        \myram/m5/dout[26] ) );
  DFFPOSX1 \myram/m5/d/d27/q_reg  ( .D(\myram/m5/mux_out[27] ), .CLK(clk), .Q(
        \myram/m5/dout[27] ) );
  DFFPOSX1 \myram/m5/d/d28/q_reg  ( .D(\myram/m5/mux_out[28] ), .CLK(clk), .Q(
        \myram/m5/dout[28] ) );
  DFFPOSX1 \myram/m5/d/d29/q_reg  ( .D(\myram/m5/mux_out[29] ), .CLK(clk), .Q(
        \myram/m5/dout[29] ) );
  DFFPOSX1 \myram/m5/d/d30/q_reg  ( .D(\myram/m5/mux_out[30] ), .CLK(clk), .Q(
        \myram/m5/dout[30] ) );
  DFFPOSX1 \myram/m5/d/d31/q_reg  ( .D(\myram/m5/mux_out[31] ), .CLK(clk), .Q(
        \myram/m5/dout[31] ) );
  DFFPOSX1 \myram/m4/d/d0/q_reg  ( .D(\myram/m4/mux_out[0] ), .CLK(clk), .Q(
        \myram/m4/dout[0] ) );
  DFFPOSX1 \myram/m4/d/d1/q_reg  ( .D(\myram/m4/mux_out[1] ), .CLK(clk), .Q(
        \myram/m4/dout[1] ) );
  DFFPOSX1 \myram/m4/d/d2/q_reg  ( .D(\myram/m4/mux_out[2] ), .CLK(clk), .Q(
        \myram/m4/dout[2] ) );
  DFFPOSX1 \myram/m4/d/d3/q_reg  ( .D(\myram/m4/mux_out[3] ), .CLK(clk), .Q(
        \myram/m4/dout[3] ) );
  DFFPOSX1 \myram/m4/d/d4/q_reg  ( .D(\myram/m4/mux_out[4] ), .CLK(clk), .Q(
        \myram/m4/dout[4] ) );
  DFFPOSX1 \myram/m4/d/d5/q_reg  ( .D(\myram/m4/mux_out[5] ), .CLK(clk), .Q(
        \myram/m4/dout[5] ) );
  DFFPOSX1 \myram/m4/d/d6/q_reg  ( .D(\myram/m4/mux_out[6] ), .CLK(clk), .Q(
        \myram/m4/dout[6] ) );
  DFFPOSX1 \myram/m4/d/d7/q_reg  ( .D(\myram/m4/mux_out[7] ), .CLK(clk), .Q(
        \myram/m4/dout[7] ) );
  DFFPOSX1 \myram/m4/d/d8/q_reg  ( .D(\myram/m4/mux_out[8] ), .CLK(clk), .Q(
        \myram/m4/dout[8] ) );
  DFFPOSX1 \myram/m4/d/d9/q_reg  ( .D(\myram/m4/mux_out[9] ), .CLK(clk), .Q(
        \myram/m4/dout[9] ) );
  DFFPOSX1 \myram/m4/d/d10/q_reg  ( .D(\myram/m4/mux_out[10] ), .CLK(clk), .Q(
        \myram/m4/dout[10] ) );
  DFFPOSX1 \myram/m4/d/d11/q_reg  ( .D(\myram/m4/mux_out[11] ), .CLK(clk), .Q(
        \myram/m4/dout[11] ) );
  DFFPOSX1 \myram/m4/d/d12/q_reg  ( .D(\myram/m4/mux_out[12] ), .CLK(clk), .Q(
        \myram/m4/dout[12] ) );
  DFFPOSX1 \myram/m4/d/d13/q_reg  ( .D(\myram/m4/mux_out[13] ), .CLK(clk), .Q(
        \myram/m4/dout[13] ) );
  DFFPOSX1 \myram/m4/d/d14/q_reg  ( .D(\myram/m4/mux_out[14] ), .CLK(clk), .Q(
        \myram/m4/dout[14] ) );
  DFFPOSX1 \myram/m4/d/d15/q_reg  ( .D(\myram/m4/mux_out[15] ), .CLK(clk), .Q(
        \myram/m4/dout[15] ) );
  DFFPOSX1 \myram/m4/d/d16/q_reg  ( .D(\myram/m4/mux_out[16] ), .CLK(clk), .Q(
        \myram/m4/dout[16] ) );
  DFFPOSX1 \myram/m4/d/d17/q_reg  ( .D(\myram/m4/mux_out[17] ), .CLK(clk), .Q(
        \myram/m4/dout[17] ) );
  DFFPOSX1 \myram/m4/d/d18/q_reg  ( .D(\myram/m4/mux_out[18] ), .CLK(clk), .Q(
        \myram/m4/dout[18] ) );
  DFFPOSX1 \myram/m4/d/d19/q_reg  ( .D(\myram/m4/mux_out[19] ), .CLK(clk), .Q(
        \myram/m4/dout[19] ) );
  DFFPOSX1 \myram/m4/d/d20/q_reg  ( .D(\myram/m4/mux_out[20] ), .CLK(clk), .Q(
        \myram/m4/dout[20] ) );
  DFFPOSX1 \myram/m4/d/d21/q_reg  ( .D(\myram/m4/mux_out[21] ), .CLK(clk), .Q(
        \myram/m4/dout[21] ) );
  DFFPOSX1 \myram/m4/d/d22/q_reg  ( .D(\myram/m4/mux_out[22] ), .CLK(clk), .Q(
        \myram/m4/dout[22] ) );
  DFFPOSX1 \myram/m4/d/d23/q_reg  ( .D(\myram/m4/mux_out[23] ), .CLK(clk), .Q(
        \myram/m4/dout[23] ) );
  DFFPOSX1 \myram/m4/d/d24/q_reg  ( .D(\myram/m4/mux_out[24] ), .CLK(clk), .Q(
        \myram/m4/dout[24] ) );
  DFFPOSX1 \myram/m4/d/d25/q_reg  ( .D(\myram/m4/mux_out[25] ), .CLK(clk), .Q(
        \myram/m4/dout[25] ) );
  DFFPOSX1 \myram/m4/d/d26/q_reg  ( .D(\myram/m4/mux_out[26] ), .CLK(clk), .Q(
        \myram/m4/dout[26] ) );
  DFFPOSX1 \myram/m4/d/d27/q_reg  ( .D(\myram/m4/mux_out[27] ), .CLK(clk), .Q(
        \myram/m4/dout[27] ) );
  DFFPOSX1 \myram/m4/d/d28/q_reg  ( .D(\myram/m4/mux_out[28] ), .CLK(clk), .Q(
        \myram/m4/dout[28] ) );
  DFFPOSX1 \myram/m4/d/d29/q_reg  ( .D(\myram/m4/mux_out[29] ), .CLK(clk), .Q(
        \myram/m4/dout[29] ) );
  DFFPOSX1 \myram/m4/d/d30/q_reg  ( .D(\myram/m4/mux_out[30] ), .CLK(clk), .Q(
        \myram/m4/dout[30] ) );
  DFFPOSX1 \myram/m4/d/d31/q_reg  ( .D(\myram/m4/mux_out[31] ), .CLK(clk), .Q(
        \myram/m4/dout[31] ) );
  DFFPOSX1 \myram/m3/d/d0/q_reg  ( .D(\myram/m3/mux_out[0] ), .CLK(clk), .Q(
        \myram/m3/dout[0] ) );
  DFFPOSX1 \myram/m3/d/d1/q_reg  ( .D(\myram/m3/mux_out[1] ), .CLK(clk), .Q(
        \myram/m3/dout[1] ) );
  DFFPOSX1 \myram/m3/d/d2/q_reg  ( .D(\myram/m3/mux_out[2] ), .CLK(clk), .Q(
        \myram/m3/dout[2] ) );
  DFFPOSX1 \myram/m3/d/d3/q_reg  ( .D(\myram/m3/mux_out[3] ), .CLK(clk), .Q(
        \myram/m3/dout[3] ) );
  DFFPOSX1 \myram/m3/d/d4/q_reg  ( .D(\myram/m3/mux_out[4] ), .CLK(clk), .Q(
        \myram/m3/dout[4] ) );
  DFFPOSX1 \myram/m3/d/d5/q_reg  ( .D(\myram/m3/mux_out[5] ), .CLK(clk), .Q(
        \myram/m3/dout[5] ) );
  DFFPOSX1 \myram/m3/d/d6/q_reg  ( .D(\myram/m3/mux_out[6] ), .CLK(clk), .Q(
        \myram/m3/dout[6] ) );
  DFFPOSX1 \myram/m3/d/d7/q_reg  ( .D(\myram/m3/mux_out[7] ), .CLK(clk), .Q(
        \myram/m3/dout[7] ) );
  DFFPOSX1 \myram/m3/d/d8/q_reg  ( .D(\myram/m3/mux_out[8] ), .CLK(clk), .Q(
        \myram/m3/dout[8] ) );
  DFFPOSX1 \myram/m3/d/d9/q_reg  ( .D(\myram/m3/mux_out[9] ), .CLK(clk), .Q(
        \myram/m3/dout[9] ) );
  DFFPOSX1 \myram/m3/d/d10/q_reg  ( .D(\myram/m3/mux_out[10] ), .CLK(clk), .Q(
        \myram/m3/dout[10] ) );
  DFFPOSX1 \myram/m3/d/d11/q_reg  ( .D(\myram/m3/mux_out[11] ), .CLK(clk), .Q(
        \myram/m3/dout[11] ) );
  DFFPOSX1 \myram/m3/d/d12/q_reg  ( .D(\myram/m3/mux_out[12] ), .CLK(clk), .Q(
        \myram/m3/dout[12] ) );
  DFFPOSX1 \myram/m3/d/d13/q_reg  ( .D(\myram/m3/mux_out[13] ), .CLK(clk), .Q(
        \myram/m3/dout[13] ) );
  DFFPOSX1 \myram/m3/d/d14/q_reg  ( .D(\myram/m3/mux_out[14] ), .CLK(clk), .Q(
        \myram/m3/dout[14] ) );
  DFFPOSX1 \myram/m3/d/d15/q_reg  ( .D(\myram/m3/mux_out[15] ), .CLK(clk), .Q(
        \myram/m3/dout[15] ) );
  DFFPOSX1 \myram/m3/d/d16/q_reg  ( .D(\myram/m3/mux_out[16] ), .CLK(clk), .Q(
        \myram/m3/dout[16] ) );
  DFFPOSX1 \myram/m3/d/d17/q_reg  ( .D(\myram/m3/mux_out[17] ), .CLK(clk), .Q(
        \myram/m3/dout[17] ) );
  DFFPOSX1 \myram/m3/d/d18/q_reg  ( .D(\myram/m3/mux_out[18] ), .CLK(clk), .Q(
        \myram/m3/dout[18] ) );
  DFFPOSX1 \myram/m3/d/d19/q_reg  ( .D(\myram/m3/mux_out[19] ), .CLK(clk), .Q(
        \myram/m3/dout[19] ) );
  DFFPOSX1 \myram/m3/d/d20/q_reg  ( .D(\myram/m3/mux_out[20] ), .CLK(clk), .Q(
        \myram/m3/dout[20] ) );
  DFFPOSX1 \myram/m3/d/d21/q_reg  ( .D(\myram/m3/mux_out[21] ), .CLK(clk), .Q(
        \myram/m3/dout[21] ) );
  DFFPOSX1 \myram/m3/d/d22/q_reg  ( .D(\myram/m3/mux_out[22] ), .CLK(clk), .Q(
        \myram/m3/dout[22] ) );
  DFFPOSX1 \myram/m3/d/d23/q_reg  ( .D(\myram/m3/mux_out[23] ), .CLK(clk), .Q(
        \myram/m3/dout[23] ) );
  DFFPOSX1 \myram/m3/d/d24/q_reg  ( .D(\myram/m3/mux_out[24] ), .CLK(clk), .Q(
        \myram/m3/dout[24] ) );
  DFFPOSX1 \myram/m3/d/d25/q_reg  ( .D(\myram/m3/mux_out[25] ), .CLK(clk), .Q(
        \myram/m3/dout[25] ) );
  DFFPOSX1 \myram/m3/d/d26/q_reg  ( .D(\myram/m3/mux_out[26] ), .CLK(clk), .Q(
        \myram/m3/dout[26] ) );
  DFFPOSX1 \myram/m3/d/d27/q_reg  ( .D(\myram/m3/mux_out[27] ), .CLK(clk), .Q(
        \myram/m3/dout[27] ) );
  DFFPOSX1 \myram/m3/d/d28/q_reg  ( .D(\myram/m3/mux_out[28] ), .CLK(clk), .Q(
        \myram/m3/dout[28] ) );
  DFFPOSX1 \myram/m3/d/d29/q_reg  ( .D(\myram/m3/mux_out[29] ), .CLK(clk), .Q(
        \myram/m3/dout[29] ) );
  DFFPOSX1 \myram/m3/d/d30/q_reg  ( .D(\myram/m3/mux_out[30] ), .CLK(clk), .Q(
        \myram/m3/dout[30] ) );
  DFFPOSX1 \myram/m3/d/d31/q_reg  ( .D(\myram/m3/mux_out[31] ), .CLK(clk), .Q(
        \myram/m3/dout[31] ) );
  DFFPOSX1 \myram/m2/d/d0/q_reg  ( .D(\myram/m2/mux_out[0] ), .CLK(clk), .Q(
        \myram/m2/dout[0] ) );
  DFFPOSX1 \myram/m2/d/d1/q_reg  ( .D(\myram/m2/mux_out[1] ), .CLK(clk), .Q(
        \myram/m2/dout[1] ) );
  DFFPOSX1 \myram/m2/d/d2/q_reg  ( .D(\myram/m2/mux_out[2] ), .CLK(clk), .Q(
        \myram/m2/dout[2] ) );
  DFFPOSX1 \myram/m2/d/d3/q_reg  ( .D(\myram/m2/mux_out[3] ), .CLK(clk), .Q(
        \myram/m2/dout[3] ) );
  DFFPOSX1 \myram/m2/d/d4/q_reg  ( .D(\myram/m2/mux_out[4] ), .CLK(clk), .Q(
        \myram/m2/dout[4] ) );
  DFFPOSX1 \myram/m2/d/d5/q_reg  ( .D(\myram/m2/mux_out[5] ), .CLK(clk), .Q(
        \myram/m2/dout[5] ) );
  DFFPOSX1 \myram/m2/d/d6/q_reg  ( .D(\myram/m2/mux_out[6] ), .CLK(clk), .Q(
        \myram/m2/dout[6] ) );
  DFFPOSX1 \myram/m2/d/d7/q_reg  ( .D(\myram/m2/mux_out[7] ), .CLK(clk), .Q(
        \myram/m2/dout[7] ) );
  DFFPOSX1 \myram/m2/d/d8/q_reg  ( .D(\myram/m2/mux_out[8] ), .CLK(clk), .Q(
        \myram/m2/dout[8] ) );
  DFFPOSX1 \myram/m2/d/d9/q_reg  ( .D(\myram/m2/mux_out[9] ), .CLK(clk), .Q(
        \myram/m2/dout[9] ) );
  DFFPOSX1 \myram/m2/d/d10/q_reg  ( .D(\myram/m2/mux_out[10] ), .CLK(clk), .Q(
        \myram/m2/dout[10] ) );
  DFFPOSX1 \myram/m2/d/d11/q_reg  ( .D(\myram/m2/mux_out[11] ), .CLK(clk), .Q(
        \myram/m2/dout[11] ) );
  DFFPOSX1 \myram/m2/d/d12/q_reg  ( .D(\myram/m2/mux_out[12] ), .CLK(clk), .Q(
        \myram/m2/dout[12] ) );
  DFFPOSX1 \myram/m2/d/d13/q_reg  ( .D(\myram/m2/mux_out[13] ), .CLK(clk), .Q(
        \myram/m2/dout[13] ) );
  DFFPOSX1 \myram/m2/d/d14/q_reg  ( .D(\myram/m2/mux_out[14] ), .CLK(clk), .Q(
        \myram/m2/dout[14] ) );
  DFFPOSX1 \myram/m2/d/d15/q_reg  ( .D(\myram/m2/mux_out[15] ), .CLK(clk), .Q(
        \myram/m2/dout[15] ) );
  DFFPOSX1 \myram/m2/d/d16/q_reg  ( .D(\myram/m2/mux_out[16] ), .CLK(clk), .Q(
        \myram/m2/dout[16] ) );
  DFFPOSX1 \myram/m2/d/d17/q_reg  ( .D(\myram/m2/mux_out[17] ), .CLK(clk), .Q(
        \myram/m2/dout[17] ) );
  DFFPOSX1 \myram/m2/d/d18/q_reg  ( .D(\myram/m2/mux_out[18] ), .CLK(clk), .Q(
        \myram/m2/dout[18] ) );
  DFFPOSX1 \myram/m2/d/d19/q_reg  ( .D(\myram/m2/mux_out[19] ), .CLK(clk), .Q(
        \myram/m2/dout[19] ) );
  DFFPOSX1 \myram/m2/d/d20/q_reg  ( .D(\myram/m2/mux_out[20] ), .CLK(clk), .Q(
        \myram/m2/dout[20] ) );
  DFFPOSX1 \myram/m2/d/d21/q_reg  ( .D(\myram/m2/mux_out[21] ), .CLK(clk), .Q(
        \myram/m2/dout[21] ) );
  DFFPOSX1 \myram/m2/d/d22/q_reg  ( .D(\myram/m2/mux_out[22] ), .CLK(clk), .Q(
        \myram/m2/dout[22] ) );
  DFFPOSX1 \myram/m2/d/d23/q_reg  ( .D(\myram/m2/mux_out[23] ), .CLK(clk), .Q(
        \myram/m2/dout[23] ) );
  DFFPOSX1 \myram/m2/d/d24/q_reg  ( .D(\myram/m2/mux_out[24] ), .CLK(clk), .Q(
        \myram/m2/dout[24] ) );
  DFFPOSX1 \myram/m2/d/d25/q_reg  ( .D(\myram/m2/mux_out[25] ), .CLK(clk), .Q(
        \myram/m2/dout[25] ) );
  DFFPOSX1 \myram/m2/d/d26/q_reg  ( .D(\myram/m2/mux_out[26] ), .CLK(clk), .Q(
        \myram/m2/dout[26] ) );
  DFFPOSX1 \myram/m2/d/d27/q_reg  ( .D(\myram/m2/mux_out[27] ), .CLK(clk), .Q(
        \myram/m2/dout[27] ) );
  DFFPOSX1 \myram/m2/d/d28/q_reg  ( .D(\myram/m2/mux_out[28] ), .CLK(clk), .Q(
        \myram/m2/dout[28] ) );
  DFFPOSX1 \myram/m2/d/d29/q_reg  ( .D(\myram/m2/mux_out[29] ), .CLK(clk), .Q(
        \myram/m2/dout[29] ) );
  DFFPOSX1 \myram/m2/d/d30/q_reg  ( .D(\myram/m2/mux_out[30] ), .CLK(clk), .Q(
        \myram/m2/dout[30] ) );
  DFFPOSX1 \myram/m2/d/d31/q_reg  ( .D(\myram/m2/mux_out[31] ), .CLK(clk), .Q(
        \myram/m2/dout[31] ) );
  DFFPOSX1 \myram/m1/d/d0/q_reg  ( .D(\myram/m1/mux_out[0] ), .CLK(clk), .Q(
        \myram/m1/dout[0] ) );
  DFFPOSX1 \myram/m1/d/d1/q_reg  ( .D(\myram/m1/mux_out[1] ), .CLK(clk), .Q(
        \myram/m1/dout[1] ) );
  DFFPOSX1 \myram/m1/d/d2/q_reg  ( .D(\myram/m1/mux_out[2] ), .CLK(clk), .Q(
        \myram/m1/dout[2] ) );
  DFFPOSX1 \myram/m1/d/d3/q_reg  ( .D(\myram/m1/mux_out[3] ), .CLK(clk), .Q(
        \myram/m1/dout[3] ) );
  DFFPOSX1 \myram/m1/d/d4/q_reg  ( .D(\myram/m1/mux_out[4] ), .CLK(clk), .Q(
        \myram/m1/dout[4] ) );
  DFFPOSX1 \myram/m1/d/d5/q_reg  ( .D(\myram/m1/mux_out[5] ), .CLK(clk), .Q(
        \myram/m1/dout[5] ) );
  DFFPOSX1 \myram/m1/d/d6/q_reg  ( .D(\myram/m1/mux_out[6] ), .CLK(clk), .Q(
        \myram/m1/dout[6] ) );
  DFFPOSX1 \myram/m1/d/d7/q_reg  ( .D(\myram/m1/mux_out[7] ), .CLK(clk), .Q(
        \myram/m1/dout[7] ) );
  DFFPOSX1 \myram/m1/d/d8/q_reg  ( .D(\myram/m1/mux_out[8] ), .CLK(clk), .Q(
        \myram/m1/dout[8] ) );
  DFFPOSX1 \myram/m1/d/d9/q_reg  ( .D(\myram/m1/mux_out[9] ), .CLK(clk), .Q(
        \myram/m1/dout[9] ) );
  DFFPOSX1 \myram/m1/d/d10/q_reg  ( .D(\myram/m1/mux_out[10] ), .CLK(clk), .Q(
        \myram/m1/dout[10] ) );
  DFFPOSX1 \myram/m1/d/d11/q_reg  ( .D(\myram/m1/mux_out[11] ), .CLK(clk), .Q(
        \myram/m1/dout[11] ) );
  DFFPOSX1 \myram/m1/d/d12/q_reg  ( .D(\myram/m1/mux_out[12] ), .CLK(clk), .Q(
        \myram/m1/dout[12] ) );
  DFFPOSX1 \myram/m1/d/d13/q_reg  ( .D(\myram/m1/mux_out[13] ), .CLK(clk), .Q(
        \myram/m1/dout[13] ) );
  DFFPOSX1 \myram/m1/d/d14/q_reg  ( .D(\myram/m1/mux_out[14] ), .CLK(clk), .Q(
        \myram/m1/dout[14] ) );
  DFFPOSX1 \myram/m1/d/d15/q_reg  ( .D(\myram/m1/mux_out[15] ), .CLK(clk), .Q(
        \myram/m1/dout[15] ) );
  DFFPOSX1 \myram/m1/d/d16/q_reg  ( .D(\myram/m1/mux_out[16] ), .CLK(clk), .Q(
        \myram/m1/dout[16] ) );
  DFFPOSX1 \myram/m1/d/d17/q_reg  ( .D(\myram/m1/mux_out[17] ), .CLK(clk), .Q(
        \myram/m1/dout[17] ) );
  DFFPOSX1 \myram/m1/d/d18/q_reg  ( .D(\myram/m1/mux_out[18] ), .CLK(clk), .Q(
        \myram/m1/dout[18] ) );
  DFFPOSX1 \myram/m1/d/d19/q_reg  ( .D(\myram/m1/mux_out[19] ), .CLK(clk), .Q(
        \myram/m1/dout[19] ) );
  DFFPOSX1 \myram/m1/d/d20/q_reg  ( .D(\myram/m1/mux_out[20] ), .CLK(clk), .Q(
        \myram/m1/dout[20] ) );
  DFFPOSX1 \myram/m1/d/d21/q_reg  ( .D(\myram/m1/mux_out[21] ), .CLK(clk), .Q(
        \myram/m1/dout[21] ) );
  DFFPOSX1 \myram/m1/d/d22/q_reg  ( .D(\myram/m1/mux_out[22] ), .CLK(clk), .Q(
        \myram/m1/dout[22] ) );
  DFFPOSX1 \myram/m1/d/d23/q_reg  ( .D(\myram/m1/mux_out[23] ), .CLK(clk), .Q(
        \myram/m1/dout[23] ) );
  DFFPOSX1 \myram/m1/d/d24/q_reg  ( .D(\myram/m1/mux_out[24] ), .CLK(clk), .Q(
        \myram/m1/dout[24] ) );
  DFFPOSX1 \myram/m1/d/d25/q_reg  ( .D(\myram/m1/mux_out[25] ), .CLK(clk), .Q(
        \myram/m1/dout[25] ) );
  DFFPOSX1 \myram/m1/d/d26/q_reg  ( .D(\myram/m1/mux_out[26] ), .CLK(clk), .Q(
        \myram/m1/dout[26] ) );
  DFFPOSX1 \myram/m1/d/d27/q_reg  ( .D(\myram/m1/mux_out[27] ), .CLK(clk), .Q(
        \myram/m1/dout[27] ) );
  DFFPOSX1 \myram/m1/d/d28/q_reg  ( .D(\myram/m1/mux_out[28] ), .CLK(clk), .Q(
        \myram/m1/dout[28] ) );
  DFFPOSX1 \myram/m1/d/d29/q_reg  ( .D(\myram/m1/mux_out[29] ), .CLK(clk), .Q(
        \myram/m1/dout[29] ) );
  DFFPOSX1 \myram/m1/d/d30/q_reg  ( .D(\myram/m1/mux_out[30] ), .CLK(clk), .Q(
        \myram/m1/dout[30] ) );
  DFFPOSX1 \myram/m1/d/d31/q_reg  ( .D(\myram/m1/mux_out[31] ), .CLK(clk), .Q(
        \myram/m1/dout[31] ) );
  NOR3X1 \myram/ds/d1/d1/U7  ( .A(n839), .B(n210), .C(n209), .Y(
        \myram/sel_s[12] ) );
  NOR3X1 \myram/ds/d1/d1/U6  ( .A(n838), .B(n210), .C(n839), .Y(
        \myram/sel_s[13] ) );
  NOR3X1 \myram/ds/d1/d1/U5  ( .A(n836), .B(n209), .C(n839), .Y(
        \myram/sel_s[14] ) );
  NOR3X1 \myram/ds/d1/d1/U4  ( .A(n836), .B(n839), .C(n838), .Y(
        \myram/sel_s[15] ) );
  NOR3X1 \myram/ds/d1/d0/U7  ( .A(n203), .B(n210), .C(n209), .Y(
        \myram/sel_s[8] ) );
  NOR3X1 \myram/ds/d1/d0/U6  ( .A(n838), .B(n210), .C(n203), .Y(
        \myram/sel_s[9] ) );
  NOR3X1 \myram/ds/d1/d0/U5  ( .A(n836), .B(n209), .C(n203), .Y(
        \myram/sel_s[10] ) );
  NOR3X1 \myram/ds/d1/d0/U4  ( .A(n836), .B(n203), .C(n838), .Y(
        \myram/sel_s[11] ) );
  NOR3X1 \myram/ds/d0/d1/U7  ( .A(n837), .B(n210), .C(n209), .Y(
        \myram/sel_s[4] ) );
  NOR3X1 \myram/ds/d0/d1/U6  ( .A(n838), .B(n210), .C(n837), .Y(
        \myram/sel_s[5] ) );
  NOR3X1 \myram/ds/d0/d1/U5  ( .A(n836), .B(n209), .C(n837), .Y(
        \myram/sel_s[6] ) );
  NOR3X1 \myram/ds/d0/d1/U4  ( .A(n836), .B(n837), .C(n838), .Y(
        \myram/sel_s[7] ) );
  NOR3X1 \myram/ds/d0/d0/U7  ( .A(n204), .B(n210), .C(n209), .Y(
        \myram/sel_s[0] ) );
  NOR3X1 \myram/ds/d0/d0/U6  ( .A(n838), .B(n210), .C(n204), .Y(
        \myram/sel_s[1] ) );
  NOR3X1 \myram/ds/d0/d0/U5  ( .A(n836), .B(n209), .C(n204), .Y(
        \myram/sel_s[2] ) );
  NOR3X1 \myram/ds/d0/d0/U4  ( .A(n836), .B(n204), .C(n838), .Y(
        \myram/sel_s[3] ) );
  NOR3X1 \myram/db/d1/d1/U7  ( .A(n835), .B(n206), .C(n205), .Y(
        \myram/sel_b[12] ) );
  NOR3X1 \myram/db/d1/d1/U6  ( .A(n833), .B(n206), .C(n835), .Y(
        \myram/sel_b[13] ) );
  NOR3X1 \myram/db/d1/d1/U5  ( .A(n832), .B(n205), .C(n835), .Y(
        \myram/sel_b[14] ) );
  NOR3X1 \myram/db/d1/d1/U4  ( .A(n832), .B(n835), .C(n833), .Y(
        \myram/sel_b[15] ) );
  NOR3X1 \myram/db/d1/d0/U7  ( .A(n194), .B(n206), .C(n205), .Y(
        \myram/sel_b[8] ) );
  NOR3X1 \myram/db/d1/d0/U6  ( .A(n833), .B(n206), .C(n194), .Y(
        \myram/sel_b[9] ) );
  NOR3X1 \myram/db/d1/d0/U5  ( .A(n832), .B(n205), .C(n194), .Y(
        \myram/sel_b[10] ) );
  NOR3X1 \myram/db/d1/d0/U4  ( .A(n832), .B(n194), .C(n833), .Y(
        \myram/sel_b[11] ) );
  NOR3X1 \myram/db/d0/d1/U7  ( .A(n834), .B(n206), .C(n205), .Y(
        \myram/sel_b[4] ) );
  NOR3X1 \myram/db/d0/d1/U6  ( .A(n833), .B(n206), .C(n834), .Y(
        \myram/sel_b[5] ) );
  NOR3X1 \myram/db/d0/d1/U5  ( .A(n832), .B(n205), .C(n834), .Y(
        \myram/sel_b[6] ) );
  NOR3X1 \myram/db/d0/d1/U4  ( .A(n832), .B(n834), .C(n833), .Y(
        \myram/sel_b[7] ) );
  NOR3X1 \myram/db/d0/d0/U7  ( .A(n205), .B(n206), .C(n193), .Y(
        \myram/sel_b[0] ) );
  NOR3X1 \myram/db/d0/d0/U6  ( .A(n833), .B(n206), .C(n193), .Y(
        \myram/sel_b[1] ) );
  NOR3X1 \myram/db/d0/d0/U5  ( .A(n832), .B(n205), .C(n193), .Y(
        \myram/sel_b[2] ) );
  NOR3X1 \myram/db/d0/d0/U4  ( .A(n832), .B(n193), .C(n833), .Y(
        \myram/sel_b[3] ) );
  NOR3X1 \myram/da/d1/d1/U7  ( .A(n831), .B(n208), .C(n207), .Y(
        \myram/sel_a[12] ) );
  NOR3X1 \myram/da/d1/d1/U6  ( .A(n829), .B(n208), .C(n831), .Y(
        \myram/sel_a[13] ) );
  NOR3X1 \myram/da/d1/d1/U5  ( .A(n828), .B(n207), .C(n831), .Y(
        \myram/sel_a[14] ) );
  NOR3X1 \myram/da/d1/d1/U4  ( .A(n828), .B(n831), .C(n829), .Y(
        \myram/sel_a[15] ) );
  NOR3X1 \myram/da/d1/d0/U7  ( .A(n191), .B(n208), .C(n207), .Y(
        \myram/sel_a[8] ) );
  NOR3X1 \myram/da/d1/d0/U6  ( .A(n829), .B(n208), .C(n191), .Y(
        \myram/sel_a[9] ) );
  NOR3X1 \myram/da/d1/d0/U5  ( .A(n828), .B(n207), .C(n191), .Y(
        \myram/sel_a[10] ) );
  NOR3X1 \myram/da/d1/d0/U4  ( .A(n828), .B(n191), .C(n829), .Y(
        \myram/sel_a[11] ) );
  NOR3X1 \myram/da/d0/d1/U7  ( .A(n830), .B(n208), .C(n207), .Y(
        \myram/sel_a[4] ) );
  NOR3X1 \myram/da/d0/d1/U6  ( .A(n829), .B(n208), .C(n830), .Y(
        \myram/sel_a[5] ) );
  NOR3X1 \myram/da/d0/d1/U5  ( .A(n828), .B(n207), .C(n830), .Y(
        \myram/sel_a[6] ) );
  NOR3X1 \myram/da/d0/d1/U4  ( .A(n828), .B(n830), .C(n829), .Y(
        \myram/sel_a[7] ) );
  TBUFX2 \myram/m15/tb/t31/b1  ( .A(n822), .EN(n245), .Y(b[31]) );
  TBUFX2 \myram/m15/tb/t30/b1  ( .A(n821), .EN(n245), .Y(b[30]) );
  TBUFX2 \myram/m15/tb/t29/b1  ( .A(n820), .EN(n245), .Y(b[29]) );
  TBUFX2 \myram/m15/tb/t28/b1  ( .A(n819), .EN(n245), .Y(b[28]) );
  TBUFX2 \myram/m15/tb/t27/b1  ( .A(n818), .EN(n245), .Y(b[27]) );
  TBUFX2 \myram/m15/tb/t26/b1  ( .A(n817), .EN(n245), .Y(b[26]) );
  TBUFX2 \myram/m15/tb/t25/b1  ( .A(n816), .EN(n245), .Y(b[25]) );
  TBUFX2 \myram/m15/tb/t24/b1  ( .A(n815), .EN(n245), .Y(b[24]) );
  TBUFX2 \myram/m15/tb/t23/b1  ( .A(n814), .EN(n245), .Y(b[23]) );
  TBUFX2 \myram/m15/tb/t22/b1  ( .A(n813), .EN(n245), .Y(b[22]) );
  TBUFX2 \myram/m15/tb/t21/b1  ( .A(n812), .EN(n245), .Y(b[21]) );
  TBUFX2 \myram/m15/tb/t20/b1  ( .A(n811), .EN(n245), .Y(b[20]) );
  TBUFX2 \myram/m15/tb/t19/b1  ( .A(n810), .EN(n245), .Y(b[19]) );
  TBUFX2 \myram/m15/tb/t18/b1  ( .A(n809), .EN(n245), .Y(b[18]) );
  TBUFX2 \myram/m15/tb/t17/b1  ( .A(n808), .EN(n245), .Y(b[17]) );
  TBUFX2 \myram/m15/tb/t16/b1  ( .A(n807), .EN(n245), .Y(b[16]) );
  TBUFX2 \myram/m15/tb/t15/b1  ( .A(n806), .EN(n245), .Y(b[15]) );
  TBUFX2 \myram/m15/tb/t14/b1  ( .A(n805), .EN(n245), .Y(b[14]) );
  TBUFX2 \myram/m15/tb/t13/b1  ( .A(n804), .EN(n245), .Y(b[13]) );
  TBUFX2 \myram/m15/tb/t12/b1  ( .A(n803), .EN(n244), .Y(b[12]) );
  TBUFX2 \myram/m15/tb/t11/b1  ( .A(n802), .EN(n244), .Y(b[11]) );
  TBUFX2 \myram/m15/tb/t10/b1  ( .A(n801), .EN(n244), .Y(b[10]) );
  TBUFX2 \myram/m15/tb/t9/b1  ( .A(n800), .EN(n244), .Y(b[9]) );
  TBUFX2 \myram/m15/tb/t8/b1  ( .A(n799), .EN(n244), .Y(b[8]) );
  TBUFX2 \myram/m15/tb/t7/b1  ( .A(n798), .EN(n244), .Y(b[7]) );
  TBUFX2 \myram/m15/tb/t6/b1  ( .A(n797), .EN(n244), .Y(b[6]) );
  TBUFX2 \myram/m15/tb/t5/b1  ( .A(n796), .EN(n244), .Y(b[5]) );
  INVX1 \myram/m15/tb/t4/U1  ( .A(\myram/m15/dout[4] ), .Y(n827) );
  TBUFX2 \myram/m15/tb/t4/b1  ( .A(n827), .EN(n244), .Y(b[4]) );
  INVX1 \myram/m15/tb/t3/U1  ( .A(\myram/m15/dout[3] ), .Y(n826) );
  TBUFX2 \myram/m15/tb/t3/b1  ( .A(n826), .EN(n244), .Y(b[3]) );
  INVX1 \myram/m15/tb/t2/U1  ( .A(\myram/m15/dout[2] ), .Y(n825) );
  TBUFX2 \myram/m15/tb/t2/b1  ( .A(n825), .EN(n244), .Y(b[2]) );
  INVX1 \myram/m15/tb/t1/U1  ( .A(\myram/m15/dout[1] ), .Y(n824) );
  TBUFX2 \myram/m15/tb/t1/b1  ( .A(n824), .EN(n244), .Y(b[1]) );
  INVX1 \myram/m15/tb/t0/U1  ( .A(\myram/m15/dout[0] ), .Y(n823) );
  TBUFX2 \myram/m15/tb/t0/b1  ( .A(n823), .EN(n244), .Y(b[0]) );
  INVX1 \myram/m15/ta/t31/U1  ( .A(\myram/m15/dout[31] ), .Y(n822) );
  TBUFX2 \myram/m15/ta/t31/b1  ( .A(n822), .EN(\myram/sel_a[15] ), .Y(a[31])
         );
  INVX1 \myram/m15/ta/t30/U1  ( .A(\myram/m15/dout[30] ), .Y(n821) );
  TBUFX2 \myram/m15/ta/t30/b1  ( .A(n821), .EN(\myram/sel_a[15] ), .Y(a[30])
         );
  INVX1 \myram/m15/ta/t29/U1  ( .A(\myram/m15/dout[29] ), .Y(n820) );
  TBUFX2 \myram/m15/ta/t29/b1  ( .A(n820), .EN(\myram/sel_a[15] ), .Y(a[29])
         );
  INVX1 \myram/m15/ta/t28/U1  ( .A(\myram/m15/dout[28] ), .Y(n819) );
  TBUFX2 \myram/m15/ta/t28/b1  ( .A(n819), .EN(\myram/sel_a[15] ), .Y(a[28])
         );
  INVX1 \myram/m15/ta/t27/U1  ( .A(\myram/m15/dout[27] ), .Y(n818) );
  TBUFX2 \myram/m15/ta/t27/b1  ( .A(n818), .EN(\myram/sel_a[15] ), .Y(a[27])
         );
  INVX1 \myram/m15/ta/t26/U1  ( .A(\myram/m15/dout[26] ), .Y(n817) );
  TBUFX2 \myram/m15/ta/t26/b1  ( .A(n817), .EN(\myram/sel_a[15] ), .Y(a[26])
         );
  INVX1 \myram/m15/ta/t25/U1  ( .A(\myram/m15/dout[25] ), .Y(n816) );
  TBUFX2 \myram/m15/ta/t25/b1  ( .A(n816), .EN(\myram/sel_a[15] ), .Y(a[25])
         );
  INVX1 \myram/m15/ta/t24/U1  ( .A(\myram/m15/dout[24] ), .Y(n815) );
  TBUFX2 \myram/m15/ta/t24/b1  ( .A(n815), .EN(\myram/sel_a[15] ), .Y(a[24])
         );
  INVX1 \myram/m15/ta/t23/U1  ( .A(\myram/m15/dout[23] ), .Y(n814) );
  TBUFX2 \myram/m15/ta/t23/b1  ( .A(n814), .EN(\myram/sel_a[15] ), .Y(a[23])
         );
  INVX1 \myram/m15/ta/t22/U1  ( .A(\myram/m15/dout[22] ), .Y(n813) );
  TBUFX2 \myram/m15/ta/t22/b1  ( .A(n813), .EN(\myram/sel_a[15] ), .Y(a[22])
         );
  INVX1 \myram/m15/ta/t21/U1  ( .A(\myram/m15/dout[21] ), .Y(n812) );
  TBUFX2 \myram/m15/ta/t21/b1  ( .A(n812), .EN(\myram/sel_a[15] ), .Y(a[21])
         );
  INVX1 \myram/m15/ta/t20/U1  ( .A(\myram/m15/dout[20] ), .Y(n811) );
  TBUFX2 \myram/m15/ta/t20/b1  ( .A(n811), .EN(\myram/sel_a[15] ), .Y(a[20])
         );
  INVX1 \myram/m15/ta/t19/U1  ( .A(\myram/m15/dout[19] ), .Y(n810) );
  TBUFX2 \myram/m15/ta/t19/b1  ( .A(n810), .EN(\myram/sel_a[15] ), .Y(a[19])
         );
  INVX1 \myram/m15/ta/t18/U1  ( .A(\myram/m15/dout[18] ), .Y(n809) );
  TBUFX2 \myram/m15/ta/t18/b1  ( .A(n809), .EN(\myram/sel_a[15] ), .Y(a[18])
         );
  INVX1 \myram/m15/ta/t17/U1  ( .A(\myram/m15/dout[17] ), .Y(n808) );
  TBUFX2 \myram/m15/ta/t17/b1  ( .A(n808), .EN(\myram/sel_a[15] ), .Y(a[17])
         );
  INVX1 \myram/m15/ta/t16/U1  ( .A(\myram/m15/dout[16] ), .Y(n807) );
  TBUFX2 \myram/m15/ta/t16/b1  ( .A(n807), .EN(\myram/sel_a[15] ), .Y(a[16])
         );
  INVX1 \myram/m15/ta/t15/U1  ( .A(\myram/m15/dout[15] ), .Y(n806) );
  TBUFX2 \myram/m15/ta/t15/b1  ( .A(n806), .EN(\myram/sel_a[15] ), .Y(a[15])
         );
  INVX1 \myram/m15/ta/t14/U1  ( .A(\myram/m15/dout[14] ), .Y(n805) );
  TBUFX2 \myram/m15/ta/t14/b1  ( .A(n805), .EN(\myram/sel_a[15] ), .Y(a[14])
         );
  INVX1 \myram/m15/ta/t13/U1  ( .A(\myram/m15/dout[13] ), .Y(n804) );
  TBUFX2 \myram/m15/ta/t13/b1  ( .A(n804), .EN(n212), .Y(a[13]) );
  INVX1 \myram/m15/ta/t12/U1  ( .A(\myram/m15/dout[12] ), .Y(n803) );
  TBUFX2 \myram/m15/ta/t12/b1  ( .A(n803), .EN(n212), .Y(a[12]) );
  INVX1 \myram/m15/ta/t11/U1  ( .A(\myram/m15/dout[11] ), .Y(n802) );
  TBUFX2 \myram/m15/ta/t11/b1  ( .A(n802), .EN(n212), .Y(a[11]) );
  INVX1 \myram/m15/ta/t10/U1  ( .A(\myram/m15/dout[10] ), .Y(n801) );
  TBUFX2 \myram/m15/ta/t10/b1  ( .A(n801), .EN(n212), .Y(a[10]) );
  INVX1 \myram/m15/ta/t9/U1  ( .A(\myram/m15/dout[9] ), .Y(n800) );
  TBUFX2 \myram/m15/ta/t9/b1  ( .A(n800), .EN(n212), .Y(a[9]) );
  INVX1 \myram/m15/ta/t8/U1  ( .A(\myram/m15/dout[8] ), .Y(n799) );
  TBUFX2 \myram/m15/ta/t8/b1  ( .A(n799), .EN(n212), .Y(a[8]) );
  INVX1 \myram/m15/ta/t7/U1  ( .A(\myram/m15/dout[7] ), .Y(n798) );
  TBUFX2 \myram/m15/ta/t7/b1  ( .A(n798), .EN(n212), .Y(a[7]) );
  INVX1 \myram/m15/ta/t6/U1  ( .A(\myram/m15/dout[6] ), .Y(n797) );
  TBUFX2 \myram/m15/ta/t6/b1  ( .A(n797), .EN(n212), .Y(a[6]) );
  INVX1 \myram/m15/ta/t5/U1  ( .A(\myram/m15/dout[5] ), .Y(n796) );
  TBUFX2 \myram/m15/ta/t5/b1  ( .A(n796), .EN(n212), .Y(a[5]) );
  TBUFX2 \myram/m15/ta/t4/b1  ( .A(n827), .EN(n212), .Y(a[4]) );
  TBUFX2 \myram/m15/ta/t3/b1  ( .A(n826), .EN(n212), .Y(a[3]) );
  TBUFX2 \myram/m15/ta/t2/b1  ( .A(n825), .EN(n212), .Y(a[2]) );
  TBUFX2 \myram/m15/ta/t1/b1  ( .A(n824), .EN(n212), .Y(a[1]) );
  TBUFX2 \myram/m15/ta/t0/b1  ( .A(n823), .EN(n212), .Y(a[0]) );
  TBUFX2 \myram/m14/tb/t31/b1  ( .A(n790), .EN(n248), .Y(b[31]) );
  TBUFX2 \myram/m14/tb/t30/b1  ( .A(n789), .EN(n248), .Y(b[30]) );
  TBUFX2 \myram/m14/tb/t29/b1  ( .A(n788), .EN(n248), .Y(b[29]) );
  TBUFX2 \myram/m14/tb/t28/b1  ( .A(n787), .EN(n248), .Y(b[28]) );
  TBUFX2 \myram/m14/tb/t27/b1  ( .A(n786), .EN(n248), .Y(b[27]) );
  TBUFX2 \myram/m14/tb/t26/b1  ( .A(n785), .EN(n248), .Y(b[26]) );
  TBUFX2 \myram/m14/tb/t25/b1  ( .A(n784), .EN(n248), .Y(b[25]) );
  TBUFX2 \myram/m14/tb/t24/b1  ( .A(n783), .EN(n248), .Y(b[24]) );
  TBUFX2 \myram/m14/tb/t23/b1  ( .A(n782), .EN(n248), .Y(b[23]) );
  TBUFX2 \myram/m14/tb/t22/b1  ( .A(n781), .EN(n248), .Y(b[22]) );
  TBUFX2 \myram/m14/tb/t21/b1  ( .A(n780), .EN(n248), .Y(b[21]) );
  TBUFX2 \myram/m14/tb/t20/b1  ( .A(n779), .EN(n248), .Y(b[20]) );
  TBUFX2 \myram/m14/tb/t19/b1  ( .A(n778), .EN(n248), .Y(b[19]) );
  TBUFX2 \myram/m14/tb/t18/b1  ( .A(n777), .EN(n248), .Y(b[18]) );
  TBUFX2 \myram/m14/tb/t17/b1  ( .A(n776), .EN(n248), .Y(b[17]) );
  TBUFX2 \myram/m14/tb/t16/b1  ( .A(n775), .EN(n248), .Y(b[16]) );
  TBUFX2 \myram/m14/tb/t15/b1  ( .A(n774), .EN(n248), .Y(b[15]) );
  TBUFX2 \myram/m14/tb/t14/b1  ( .A(n773), .EN(n248), .Y(b[14]) );
  TBUFX2 \myram/m14/tb/t13/b1  ( .A(n772), .EN(n248), .Y(b[13]) );
  TBUFX2 \myram/m14/tb/t12/b1  ( .A(n771), .EN(n247), .Y(b[12]) );
  TBUFX2 \myram/m14/tb/t11/b1  ( .A(n770), .EN(n247), .Y(b[11]) );
  TBUFX2 \myram/m14/tb/t10/b1  ( .A(n769), .EN(n247), .Y(b[10]) );
  TBUFX2 \myram/m14/tb/t9/b1  ( .A(n768), .EN(n247), .Y(b[9]) );
  TBUFX2 \myram/m14/tb/t8/b1  ( .A(n767), .EN(n247), .Y(b[8]) );
  TBUFX2 \myram/m14/tb/t7/b1  ( .A(n766), .EN(n247), .Y(b[7]) );
  TBUFX2 \myram/m14/tb/t6/b1  ( .A(n765), .EN(n247), .Y(b[6]) );
  TBUFX2 \myram/m14/tb/t5/b1  ( .A(n764), .EN(n247), .Y(b[5]) );
  INVX1 \myram/m14/tb/t4/U1  ( .A(\myram/m14/dout[4] ), .Y(n795) );
  TBUFX2 \myram/m14/tb/t4/b1  ( .A(n795), .EN(n247), .Y(b[4]) );
  INVX1 \myram/m14/tb/t3/U1  ( .A(\myram/m14/dout[3] ), .Y(n794) );
  TBUFX2 \myram/m14/tb/t3/b1  ( .A(n794), .EN(n247), .Y(b[3]) );
  INVX1 \myram/m14/tb/t2/U1  ( .A(\myram/m14/dout[2] ), .Y(n793) );
  TBUFX2 \myram/m14/tb/t2/b1  ( .A(n793), .EN(n247), .Y(b[2]) );
  INVX1 \myram/m14/tb/t1/U1  ( .A(\myram/m14/dout[1] ), .Y(n792) );
  TBUFX2 \myram/m14/tb/t1/b1  ( .A(n792), .EN(n247), .Y(b[1]) );
  INVX1 \myram/m14/tb/t0/U1  ( .A(\myram/m14/dout[0] ), .Y(n791) );
  TBUFX2 \myram/m14/tb/t0/b1  ( .A(n791), .EN(n247), .Y(b[0]) );
  INVX1 \myram/m14/ta/t31/U1  ( .A(\myram/m14/dout[31] ), .Y(n790) );
  TBUFX2 \myram/m14/ta/t31/b1  ( .A(n790), .EN(\myram/sel_a[14] ), .Y(a[31])
         );
  INVX1 \myram/m14/ta/t30/U1  ( .A(\myram/m14/dout[30] ), .Y(n789) );
  TBUFX2 \myram/m14/ta/t30/b1  ( .A(n789), .EN(\myram/sel_a[14] ), .Y(a[30])
         );
  INVX1 \myram/m14/ta/t29/U1  ( .A(\myram/m14/dout[29] ), .Y(n788) );
  TBUFX2 \myram/m14/ta/t29/b1  ( .A(n788), .EN(\myram/sel_a[14] ), .Y(a[29])
         );
  INVX1 \myram/m14/ta/t28/U1  ( .A(\myram/m14/dout[28] ), .Y(n787) );
  TBUFX2 \myram/m14/ta/t28/b1  ( .A(n787), .EN(\myram/sel_a[14] ), .Y(a[28])
         );
  INVX1 \myram/m14/ta/t27/U1  ( .A(\myram/m14/dout[27] ), .Y(n786) );
  TBUFX2 \myram/m14/ta/t27/b1  ( .A(n786), .EN(\myram/sel_a[14] ), .Y(a[27])
         );
  INVX1 \myram/m14/ta/t26/U1  ( .A(\myram/m14/dout[26] ), .Y(n785) );
  TBUFX2 \myram/m14/ta/t26/b1  ( .A(n785), .EN(\myram/sel_a[14] ), .Y(a[26])
         );
  INVX1 \myram/m14/ta/t25/U1  ( .A(\myram/m14/dout[25] ), .Y(n784) );
  TBUFX2 \myram/m14/ta/t25/b1  ( .A(n784), .EN(\myram/sel_a[14] ), .Y(a[25])
         );
  INVX1 \myram/m14/ta/t24/U1  ( .A(\myram/m14/dout[24] ), .Y(n783) );
  TBUFX2 \myram/m14/ta/t24/b1  ( .A(n783), .EN(\myram/sel_a[14] ), .Y(a[24])
         );
  INVX1 \myram/m14/ta/t23/U1  ( .A(\myram/m14/dout[23] ), .Y(n782) );
  TBUFX2 \myram/m14/ta/t23/b1  ( .A(n782), .EN(\myram/sel_a[14] ), .Y(a[23])
         );
  INVX1 \myram/m14/ta/t22/U1  ( .A(\myram/m14/dout[22] ), .Y(n781) );
  TBUFX2 \myram/m14/ta/t22/b1  ( .A(n781), .EN(\myram/sel_a[14] ), .Y(a[22])
         );
  INVX1 \myram/m14/ta/t21/U1  ( .A(\myram/m14/dout[21] ), .Y(n780) );
  TBUFX2 \myram/m14/ta/t21/b1  ( .A(n780), .EN(\myram/sel_a[14] ), .Y(a[21])
         );
  INVX1 \myram/m14/ta/t20/U1  ( .A(\myram/m14/dout[20] ), .Y(n779) );
  TBUFX2 \myram/m14/ta/t20/b1  ( .A(n779), .EN(\myram/sel_a[14] ), .Y(a[20])
         );
  INVX1 \myram/m14/ta/t19/U1  ( .A(\myram/m14/dout[19] ), .Y(n778) );
  TBUFX2 \myram/m14/ta/t19/b1  ( .A(n778), .EN(\myram/sel_a[14] ), .Y(a[19])
         );
  INVX1 \myram/m14/ta/t18/U1  ( .A(\myram/m14/dout[18] ), .Y(n777) );
  TBUFX2 \myram/m14/ta/t18/b1  ( .A(n777), .EN(\myram/sel_a[14] ), .Y(a[18])
         );
  INVX1 \myram/m14/ta/t17/U1  ( .A(\myram/m14/dout[17] ), .Y(n776) );
  TBUFX2 \myram/m14/ta/t17/b1  ( .A(n776), .EN(\myram/sel_a[14] ), .Y(a[17])
         );
  INVX1 \myram/m14/ta/t16/U1  ( .A(\myram/m14/dout[16] ), .Y(n775) );
  TBUFX2 \myram/m14/ta/t16/b1  ( .A(n775), .EN(\myram/sel_a[14] ), .Y(a[16])
         );
  INVX1 \myram/m14/ta/t15/U1  ( .A(\myram/m14/dout[15] ), .Y(n774) );
  TBUFX2 \myram/m14/ta/t15/b1  ( .A(n774), .EN(\myram/sel_a[14] ), .Y(a[15])
         );
  INVX1 \myram/m14/ta/t14/U1  ( .A(\myram/m14/dout[14] ), .Y(n773) );
  TBUFX2 \myram/m14/ta/t14/b1  ( .A(n773), .EN(\myram/sel_a[14] ), .Y(a[14])
         );
  INVX1 \myram/m14/ta/t13/U1  ( .A(\myram/m14/dout[13] ), .Y(n772) );
  TBUFX2 \myram/m14/ta/t13/b1  ( .A(n772), .EN(n214), .Y(a[13]) );
  INVX1 \myram/m14/ta/t12/U1  ( .A(\myram/m14/dout[12] ), .Y(n771) );
  TBUFX2 \myram/m14/ta/t12/b1  ( .A(n771), .EN(n214), .Y(a[12]) );
  INVX1 \myram/m14/ta/t11/U1  ( .A(\myram/m14/dout[11] ), .Y(n770) );
  TBUFX2 \myram/m14/ta/t11/b1  ( .A(n770), .EN(n214), .Y(a[11]) );
  INVX1 \myram/m14/ta/t10/U1  ( .A(\myram/m14/dout[10] ), .Y(n769) );
  TBUFX2 \myram/m14/ta/t10/b1  ( .A(n769), .EN(n214), .Y(a[10]) );
  INVX1 \myram/m14/ta/t9/U1  ( .A(\myram/m14/dout[9] ), .Y(n768) );
  TBUFX2 \myram/m14/ta/t9/b1  ( .A(n768), .EN(n214), .Y(a[9]) );
  INVX1 \myram/m14/ta/t8/U1  ( .A(\myram/m14/dout[8] ), .Y(n767) );
  TBUFX2 \myram/m14/ta/t8/b1  ( .A(n767), .EN(n214), .Y(a[8]) );
  INVX1 \myram/m14/ta/t7/U1  ( .A(\myram/m14/dout[7] ), .Y(n766) );
  TBUFX2 \myram/m14/ta/t7/b1  ( .A(n766), .EN(n214), .Y(a[7]) );
  INVX1 \myram/m14/ta/t6/U1  ( .A(\myram/m14/dout[6] ), .Y(n765) );
  TBUFX2 \myram/m14/ta/t6/b1  ( .A(n765), .EN(n214), .Y(a[6]) );
  INVX1 \myram/m14/ta/t5/U1  ( .A(\myram/m14/dout[5] ), .Y(n764) );
  TBUFX2 \myram/m14/ta/t5/b1  ( .A(n764), .EN(n214), .Y(a[5]) );
  TBUFX2 \myram/m14/ta/t4/b1  ( .A(n795), .EN(n214), .Y(a[4]) );
  TBUFX2 \myram/m14/ta/t3/b1  ( .A(n794), .EN(n214), .Y(a[3]) );
  TBUFX2 \myram/m14/ta/t2/b1  ( .A(n793), .EN(n214), .Y(a[2]) );
  TBUFX2 \myram/m14/ta/t1/b1  ( .A(n792), .EN(n214), .Y(a[1]) );
  TBUFX2 \myram/m14/ta/t0/b1  ( .A(n791), .EN(n214), .Y(a[0]) );
  TBUFX2 \myram/m13/tb/t31/b1  ( .A(n758), .EN(n251), .Y(b[31]) );
  TBUFX2 \myram/m13/tb/t30/b1  ( .A(n757), .EN(n251), .Y(b[30]) );
  TBUFX2 \myram/m13/tb/t29/b1  ( .A(n756), .EN(n251), .Y(b[29]) );
  TBUFX2 \myram/m13/tb/t28/b1  ( .A(n755), .EN(n251), .Y(b[28]) );
  TBUFX2 \myram/m13/tb/t27/b1  ( .A(n754), .EN(n251), .Y(b[27]) );
  TBUFX2 \myram/m13/tb/t26/b1  ( .A(n753), .EN(n251), .Y(b[26]) );
  TBUFX2 \myram/m13/tb/t25/b1  ( .A(n752), .EN(n251), .Y(b[25]) );
  TBUFX2 \myram/m13/tb/t24/b1  ( .A(n751), .EN(n251), .Y(b[24]) );
  TBUFX2 \myram/m13/tb/t23/b1  ( .A(n750), .EN(n251), .Y(b[23]) );
  TBUFX2 \myram/m13/tb/t22/b1  ( .A(n749), .EN(n251), .Y(b[22]) );
  TBUFX2 \myram/m13/tb/t21/b1  ( .A(n748), .EN(n251), .Y(b[21]) );
  TBUFX2 \myram/m13/tb/t20/b1  ( .A(n747), .EN(n251), .Y(b[20]) );
  TBUFX2 \myram/m13/tb/t19/b1  ( .A(n746), .EN(n251), .Y(b[19]) );
  TBUFX2 \myram/m13/tb/t18/b1  ( .A(n745), .EN(n251), .Y(b[18]) );
  TBUFX2 \myram/m13/tb/t17/b1  ( .A(n744), .EN(n251), .Y(b[17]) );
  TBUFX2 \myram/m13/tb/t16/b1  ( .A(n743), .EN(n251), .Y(b[16]) );
  TBUFX2 \myram/m13/tb/t15/b1  ( .A(n742), .EN(n251), .Y(b[15]) );
  TBUFX2 \myram/m13/tb/t14/b1  ( .A(n741), .EN(n251), .Y(b[14]) );
  TBUFX2 \myram/m13/tb/t13/b1  ( .A(n740), .EN(n251), .Y(b[13]) );
  TBUFX2 \myram/m13/tb/t12/b1  ( .A(n739), .EN(n250), .Y(b[12]) );
  TBUFX2 \myram/m13/tb/t11/b1  ( .A(n738), .EN(n250), .Y(b[11]) );
  TBUFX2 \myram/m13/tb/t10/b1  ( .A(n737), .EN(n250), .Y(b[10]) );
  TBUFX2 \myram/m13/tb/t9/b1  ( .A(n736), .EN(n250), .Y(b[9]) );
  TBUFX2 \myram/m13/tb/t8/b1  ( .A(n735), .EN(n250), .Y(b[8]) );
  TBUFX2 \myram/m13/tb/t7/b1  ( .A(n734), .EN(n250), .Y(b[7]) );
  TBUFX2 \myram/m13/tb/t6/b1  ( .A(n733), .EN(n250), .Y(b[6]) );
  TBUFX2 \myram/m13/tb/t5/b1  ( .A(n732), .EN(n250), .Y(b[5]) );
  INVX1 \myram/m13/tb/t4/U1  ( .A(\myram/m13/dout[4] ), .Y(n763) );
  TBUFX2 \myram/m13/tb/t4/b1  ( .A(n763), .EN(n250), .Y(b[4]) );
  INVX1 \myram/m13/tb/t3/U1  ( .A(\myram/m13/dout[3] ), .Y(n762) );
  TBUFX2 \myram/m13/tb/t3/b1  ( .A(n762), .EN(n250), .Y(b[3]) );
  INVX1 \myram/m13/tb/t2/U1  ( .A(\myram/m13/dout[2] ), .Y(n761) );
  TBUFX2 \myram/m13/tb/t2/b1  ( .A(n761), .EN(n250), .Y(b[2]) );
  INVX1 \myram/m13/tb/t1/U1  ( .A(\myram/m13/dout[1] ), .Y(n760) );
  TBUFX2 \myram/m13/tb/t1/b1  ( .A(n760), .EN(n250), .Y(b[1]) );
  INVX1 \myram/m13/tb/t0/U1  ( .A(\myram/m13/dout[0] ), .Y(n759) );
  TBUFX2 \myram/m13/tb/t0/b1  ( .A(n759), .EN(n250), .Y(b[0]) );
  INVX1 \myram/m13/ta/t31/U1  ( .A(\myram/m13/dout[31] ), .Y(n758) );
  TBUFX2 \myram/m13/ta/t31/b1  ( .A(n758), .EN(\myram/sel_a[13] ), .Y(a[31])
         );
  INVX1 \myram/m13/ta/t30/U1  ( .A(\myram/m13/dout[30] ), .Y(n757) );
  TBUFX2 \myram/m13/ta/t30/b1  ( .A(n757), .EN(\myram/sel_a[13] ), .Y(a[30])
         );
  INVX1 \myram/m13/ta/t29/U1  ( .A(\myram/m13/dout[29] ), .Y(n756) );
  TBUFX2 \myram/m13/ta/t29/b1  ( .A(n756), .EN(\myram/sel_a[13] ), .Y(a[29])
         );
  INVX1 \myram/m13/ta/t28/U1  ( .A(\myram/m13/dout[28] ), .Y(n755) );
  TBUFX2 \myram/m13/ta/t28/b1  ( .A(n755), .EN(\myram/sel_a[13] ), .Y(a[28])
         );
  INVX1 \myram/m13/ta/t27/U1  ( .A(\myram/m13/dout[27] ), .Y(n754) );
  TBUFX2 \myram/m13/ta/t27/b1  ( .A(n754), .EN(\myram/sel_a[13] ), .Y(a[27])
         );
  INVX1 \myram/m13/ta/t26/U1  ( .A(\myram/m13/dout[26] ), .Y(n753) );
  TBUFX2 \myram/m13/ta/t26/b1  ( .A(n753), .EN(\myram/sel_a[13] ), .Y(a[26])
         );
  INVX1 \myram/m13/ta/t25/U1  ( .A(\myram/m13/dout[25] ), .Y(n752) );
  TBUFX2 \myram/m13/ta/t25/b1  ( .A(n752), .EN(\myram/sel_a[13] ), .Y(a[25])
         );
  INVX1 \myram/m13/ta/t24/U1  ( .A(\myram/m13/dout[24] ), .Y(n751) );
  TBUFX2 \myram/m13/ta/t24/b1  ( .A(n751), .EN(\myram/sel_a[13] ), .Y(a[24])
         );
  INVX1 \myram/m13/ta/t23/U1  ( .A(\myram/m13/dout[23] ), .Y(n750) );
  TBUFX2 \myram/m13/ta/t23/b1  ( .A(n750), .EN(\myram/sel_a[13] ), .Y(a[23])
         );
  INVX1 \myram/m13/ta/t22/U1  ( .A(\myram/m13/dout[22] ), .Y(n749) );
  TBUFX2 \myram/m13/ta/t22/b1  ( .A(n749), .EN(\myram/sel_a[13] ), .Y(a[22])
         );
  INVX1 \myram/m13/ta/t21/U1  ( .A(\myram/m13/dout[21] ), .Y(n748) );
  TBUFX2 \myram/m13/ta/t21/b1  ( .A(n748), .EN(\myram/sel_a[13] ), .Y(a[21])
         );
  INVX1 \myram/m13/ta/t20/U1  ( .A(\myram/m13/dout[20] ), .Y(n747) );
  TBUFX2 \myram/m13/ta/t20/b1  ( .A(n747), .EN(\myram/sel_a[13] ), .Y(a[20])
         );
  INVX1 \myram/m13/ta/t19/U1  ( .A(\myram/m13/dout[19] ), .Y(n746) );
  TBUFX2 \myram/m13/ta/t19/b1  ( .A(n746), .EN(\myram/sel_a[13] ), .Y(a[19])
         );
  INVX1 \myram/m13/ta/t18/U1  ( .A(\myram/m13/dout[18] ), .Y(n745) );
  TBUFX2 \myram/m13/ta/t18/b1  ( .A(n745), .EN(\myram/sel_a[13] ), .Y(a[18])
         );
  INVX1 \myram/m13/ta/t17/U1  ( .A(\myram/m13/dout[17] ), .Y(n744) );
  TBUFX2 \myram/m13/ta/t17/b1  ( .A(n744), .EN(\myram/sel_a[13] ), .Y(a[17])
         );
  INVX1 \myram/m13/ta/t16/U1  ( .A(\myram/m13/dout[16] ), .Y(n743) );
  TBUFX2 \myram/m13/ta/t16/b1  ( .A(n743), .EN(\myram/sel_a[13] ), .Y(a[16])
         );
  INVX1 \myram/m13/ta/t15/U1  ( .A(\myram/m13/dout[15] ), .Y(n742) );
  TBUFX2 \myram/m13/ta/t15/b1  ( .A(n742), .EN(\myram/sel_a[13] ), .Y(a[15])
         );
  INVX1 \myram/m13/ta/t14/U1  ( .A(\myram/m13/dout[14] ), .Y(n741) );
  TBUFX2 \myram/m13/ta/t14/b1  ( .A(n741), .EN(\myram/sel_a[13] ), .Y(a[14])
         );
  INVX1 \myram/m13/ta/t13/U1  ( .A(\myram/m13/dout[13] ), .Y(n740) );
  TBUFX2 \myram/m13/ta/t13/b1  ( .A(n740), .EN(n216), .Y(a[13]) );
  INVX1 \myram/m13/ta/t12/U1  ( .A(\myram/m13/dout[12] ), .Y(n739) );
  TBUFX2 \myram/m13/ta/t12/b1  ( .A(n739), .EN(n216), .Y(a[12]) );
  INVX1 \myram/m13/ta/t11/U1  ( .A(\myram/m13/dout[11] ), .Y(n738) );
  TBUFX2 \myram/m13/ta/t11/b1  ( .A(n738), .EN(n216), .Y(a[11]) );
  INVX1 \myram/m13/ta/t10/U1  ( .A(\myram/m13/dout[10] ), .Y(n737) );
  TBUFX2 \myram/m13/ta/t10/b1  ( .A(n737), .EN(n216), .Y(a[10]) );
  INVX1 \myram/m13/ta/t9/U1  ( .A(\myram/m13/dout[9] ), .Y(n736) );
  TBUFX2 \myram/m13/ta/t9/b1  ( .A(n736), .EN(n216), .Y(a[9]) );
  INVX1 \myram/m13/ta/t8/U1  ( .A(\myram/m13/dout[8] ), .Y(n735) );
  TBUFX2 \myram/m13/ta/t8/b1  ( .A(n735), .EN(n216), .Y(a[8]) );
  INVX1 \myram/m13/ta/t7/U1  ( .A(\myram/m13/dout[7] ), .Y(n734) );
  TBUFX2 \myram/m13/ta/t7/b1  ( .A(n734), .EN(n216), .Y(a[7]) );
  INVX1 \myram/m13/ta/t6/U1  ( .A(\myram/m13/dout[6] ), .Y(n733) );
  TBUFX2 \myram/m13/ta/t6/b1  ( .A(n733), .EN(n216), .Y(a[6]) );
  INVX1 \myram/m13/ta/t5/U1  ( .A(\myram/m13/dout[5] ), .Y(n732) );
  TBUFX2 \myram/m13/ta/t5/b1  ( .A(n732), .EN(n216), .Y(a[5]) );
  TBUFX2 \myram/m13/ta/t4/b1  ( .A(n763), .EN(n216), .Y(a[4]) );
  TBUFX2 \myram/m13/ta/t3/b1  ( .A(n762), .EN(n216), .Y(a[3]) );
  TBUFX2 \myram/m13/ta/t2/b1  ( .A(n761), .EN(n216), .Y(a[2]) );
  TBUFX2 \myram/m13/ta/t1/b1  ( .A(n760), .EN(n216), .Y(a[1]) );
  TBUFX2 \myram/m13/ta/t0/b1  ( .A(n759), .EN(n216), .Y(a[0]) );
  TBUFX2 \myram/m12/tb/t31/b1  ( .A(n726), .EN(n254), .Y(b[31]) );
  TBUFX2 \myram/m12/tb/t30/b1  ( .A(n725), .EN(n254), .Y(b[30]) );
  TBUFX2 \myram/m12/tb/t29/b1  ( .A(n724), .EN(n254), .Y(b[29]) );
  TBUFX2 \myram/m12/tb/t28/b1  ( .A(n723), .EN(n254), .Y(b[28]) );
  TBUFX2 \myram/m12/tb/t27/b1  ( .A(n722), .EN(n254), .Y(b[27]) );
  TBUFX2 \myram/m12/tb/t26/b1  ( .A(n721), .EN(n254), .Y(b[26]) );
  TBUFX2 \myram/m12/tb/t25/b1  ( .A(n720), .EN(n254), .Y(b[25]) );
  TBUFX2 \myram/m12/tb/t24/b1  ( .A(n719), .EN(n254), .Y(b[24]) );
  TBUFX2 \myram/m12/tb/t23/b1  ( .A(n718), .EN(n254), .Y(b[23]) );
  TBUFX2 \myram/m12/tb/t22/b1  ( .A(n717), .EN(n254), .Y(b[22]) );
  TBUFX2 \myram/m12/tb/t21/b1  ( .A(n716), .EN(n254), .Y(b[21]) );
  TBUFX2 \myram/m12/tb/t20/b1  ( .A(n715), .EN(n254), .Y(b[20]) );
  TBUFX2 \myram/m12/tb/t19/b1  ( .A(n714), .EN(n254), .Y(b[19]) );
  TBUFX2 \myram/m12/tb/t18/b1  ( .A(n713), .EN(n254), .Y(b[18]) );
  TBUFX2 \myram/m12/tb/t17/b1  ( .A(n712), .EN(n254), .Y(b[17]) );
  TBUFX2 \myram/m12/tb/t16/b1  ( .A(n711), .EN(n254), .Y(b[16]) );
  TBUFX2 \myram/m12/tb/t15/b1  ( .A(n710), .EN(n254), .Y(b[15]) );
  TBUFX2 \myram/m12/tb/t14/b1  ( .A(n709), .EN(n254), .Y(b[14]) );
  TBUFX2 \myram/m12/tb/t13/b1  ( .A(n708), .EN(n254), .Y(b[13]) );
  TBUFX2 \myram/m12/tb/t12/b1  ( .A(n707), .EN(n253), .Y(b[12]) );
  TBUFX2 \myram/m12/tb/t11/b1  ( .A(n706), .EN(n253), .Y(b[11]) );
  TBUFX2 \myram/m12/tb/t10/b1  ( .A(n705), .EN(n253), .Y(b[10]) );
  TBUFX2 \myram/m12/tb/t9/b1  ( .A(n704), .EN(n253), .Y(b[9]) );
  TBUFX2 \myram/m12/tb/t8/b1  ( .A(n703), .EN(n253), .Y(b[8]) );
  TBUFX2 \myram/m12/tb/t7/b1  ( .A(n702), .EN(n253), .Y(b[7]) );
  TBUFX2 \myram/m12/tb/t6/b1  ( .A(n701), .EN(n253), .Y(b[6]) );
  TBUFX2 \myram/m12/tb/t5/b1  ( .A(n700), .EN(n253), .Y(b[5]) );
  INVX1 \myram/m12/tb/t4/U1  ( .A(\myram/m12/dout[4] ), .Y(n731) );
  TBUFX2 \myram/m12/tb/t4/b1  ( .A(n731), .EN(n253), .Y(b[4]) );
  INVX1 \myram/m12/tb/t3/U1  ( .A(\myram/m12/dout[3] ), .Y(n730) );
  TBUFX2 \myram/m12/tb/t3/b1  ( .A(n730), .EN(n253), .Y(b[3]) );
  INVX1 \myram/m12/tb/t2/U1  ( .A(\myram/m12/dout[2] ), .Y(n729) );
  TBUFX2 \myram/m12/tb/t2/b1  ( .A(n729), .EN(n253), .Y(b[2]) );
  INVX1 \myram/m12/tb/t1/U1  ( .A(\myram/m12/dout[1] ), .Y(n728) );
  TBUFX2 \myram/m12/tb/t1/b1  ( .A(n728), .EN(n253), .Y(b[1]) );
  INVX1 \myram/m12/tb/t0/U1  ( .A(\myram/m12/dout[0] ), .Y(n727) );
  TBUFX2 \myram/m12/tb/t0/b1  ( .A(n727), .EN(n253), .Y(b[0]) );
  INVX1 \myram/m12/ta/t31/U1  ( .A(\myram/m12/dout[31] ), .Y(n726) );
  TBUFX2 \myram/m12/ta/t31/b1  ( .A(n726), .EN(\myram/sel_a[12] ), .Y(a[31])
         );
  INVX1 \myram/m12/ta/t30/U1  ( .A(\myram/m12/dout[30] ), .Y(n725) );
  TBUFX2 \myram/m12/ta/t30/b1  ( .A(n725), .EN(\myram/sel_a[12] ), .Y(a[30])
         );
  INVX1 \myram/m12/ta/t29/U1  ( .A(\myram/m12/dout[29] ), .Y(n724) );
  TBUFX2 \myram/m12/ta/t29/b1  ( .A(n724), .EN(\myram/sel_a[12] ), .Y(a[29])
         );
  INVX1 \myram/m12/ta/t28/U1  ( .A(\myram/m12/dout[28] ), .Y(n723) );
  TBUFX2 \myram/m12/ta/t28/b1  ( .A(n723), .EN(\myram/sel_a[12] ), .Y(a[28])
         );
  INVX1 \myram/m12/ta/t27/U1  ( .A(\myram/m12/dout[27] ), .Y(n722) );
  TBUFX2 \myram/m12/ta/t27/b1  ( .A(n722), .EN(\myram/sel_a[12] ), .Y(a[27])
         );
  INVX1 \myram/m12/ta/t26/U1  ( .A(\myram/m12/dout[26] ), .Y(n721) );
  TBUFX2 \myram/m12/ta/t26/b1  ( .A(n721), .EN(\myram/sel_a[12] ), .Y(a[26])
         );
  INVX1 \myram/m12/ta/t25/U1  ( .A(\myram/m12/dout[25] ), .Y(n720) );
  TBUFX2 \myram/m12/ta/t25/b1  ( .A(n720), .EN(\myram/sel_a[12] ), .Y(a[25])
         );
  INVX1 \myram/m12/ta/t24/U1  ( .A(\myram/m12/dout[24] ), .Y(n719) );
  TBUFX2 \myram/m12/ta/t24/b1  ( .A(n719), .EN(\myram/sel_a[12] ), .Y(a[24])
         );
  INVX1 \myram/m12/ta/t23/U1  ( .A(\myram/m12/dout[23] ), .Y(n718) );
  TBUFX2 \myram/m12/ta/t23/b1  ( .A(n718), .EN(\myram/sel_a[12] ), .Y(a[23])
         );
  INVX1 \myram/m12/ta/t22/U1  ( .A(\myram/m12/dout[22] ), .Y(n717) );
  TBUFX2 \myram/m12/ta/t22/b1  ( .A(n717), .EN(\myram/sel_a[12] ), .Y(a[22])
         );
  INVX1 \myram/m12/ta/t21/U1  ( .A(\myram/m12/dout[21] ), .Y(n716) );
  TBUFX2 \myram/m12/ta/t21/b1  ( .A(n716), .EN(\myram/sel_a[12] ), .Y(a[21])
         );
  INVX1 \myram/m12/ta/t20/U1  ( .A(\myram/m12/dout[20] ), .Y(n715) );
  TBUFX2 \myram/m12/ta/t20/b1  ( .A(n715), .EN(\myram/sel_a[12] ), .Y(a[20])
         );
  INVX1 \myram/m12/ta/t19/U1  ( .A(\myram/m12/dout[19] ), .Y(n714) );
  TBUFX2 \myram/m12/ta/t19/b1  ( .A(n714), .EN(\myram/sel_a[12] ), .Y(a[19])
         );
  INVX1 \myram/m12/ta/t18/U1  ( .A(\myram/m12/dout[18] ), .Y(n713) );
  TBUFX2 \myram/m12/ta/t18/b1  ( .A(n713), .EN(\myram/sel_a[12] ), .Y(a[18])
         );
  INVX1 \myram/m12/ta/t17/U1  ( .A(\myram/m12/dout[17] ), .Y(n712) );
  TBUFX2 \myram/m12/ta/t17/b1  ( .A(n712), .EN(\myram/sel_a[12] ), .Y(a[17])
         );
  INVX1 \myram/m12/ta/t16/U1  ( .A(\myram/m12/dout[16] ), .Y(n711) );
  TBUFX2 \myram/m12/ta/t16/b1  ( .A(n711), .EN(\myram/sel_a[12] ), .Y(a[16])
         );
  INVX1 \myram/m12/ta/t15/U1  ( .A(\myram/m12/dout[15] ), .Y(n710) );
  TBUFX2 \myram/m12/ta/t15/b1  ( .A(n710), .EN(\myram/sel_a[12] ), .Y(a[15])
         );
  INVX1 \myram/m12/ta/t14/U1  ( .A(\myram/m12/dout[14] ), .Y(n709) );
  TBUFX2 \myram/m12/ta/t14/b1  ( .A(n709), .EN(\myram/sel_a[12] ), .Y(a[14])
         );
  INVX1 \myram/m12/ta/t13/U1  ( .A(\myram/m12/dout[13] ), .Y(n708) );
  TBUFX2 \myram/m12/ta/t13/b1  ( .A(n708), .EN(n218), .Y(a[13]) );
  INVX1 \myram/m12/ta/t12/U1  ( .A(\myram/m12/dout[12] ), .Y(n707) );
  TBUFX2 \myram/m12/ta/t12/b1  ( .A(n707), .EN(n218), .Y(a[12]) );
  INVX1 \myram/m12/ta/t11/U1  ( .A(\myram/m12/dout[11] ), .Y(n706) );
  TBUFX2 \myram/m12/ta/t11/b1  ( .A(n706), .EN(n218), .Y(a[11]) );
  INVX1 \myram/m12/ta/t10/U1  ( .A(\myram/m12/dout[10] ), .Y(n705) );
  TBUFX2 \myram/m12/ta/t10/b1  ( .A(n705), .EN(n218), .Y(a[10]) );
  INVX1 \myram/m12/ta/t9/U1  ( .A(\myram/m12/dout[9] ), .Y(n704) );
  TBUFX2 \myram/m12/ta/t9/b1  ( .A(n704), .EN(n218), .Y(a[9]) );
  INVX1 \myram/m12/ta/t8/U1  ( .A(\myram/m12/dout[8] ), .Y(n703) );
  TBUFX2 \myram/m12/ta/t8/b1  ( .A(n703), .EN(n218), .Y(a[8]) );
  INVX1 \myram/m12/ta/t7/U1  ( .A(\myram/m12/dout[7] ), .Y(n702) );
  TBUFX2 \myram/m12/ta/t7/b1  ( .A(n702), .EN(n218), .Y(a[7]) );
  INVX1 \myram/m12/ta/t6/U1  ( .A(\myram/m12/dout[6] ), .Y(n701) );
  TBUFX2 \myram/m12/ta/t6/b1  ( .A(n701), .EN(n218), .Y(a[6]) );
  INVX1 \myram/m12/ta/t5/U1  ( .A(\myram/m12/dout[5] ), .Y(n700) );
  TBUFX2 \myram/m12/ta/t5/b1  ( .A(n700), .EN(n218), .Y(a[5]) );
  TBUFX2 \myram/m12/ta/t4/b1  ( .A(n731), .EN(n218), .Y(a[4]) );
  TBUFX2 \myram/m12/ta/t3/b1  ( .A(n730), .EN(n218), .Y(a[3]) );
  TBUFX2 \myram/m12/ta/t2/b1  ( .A(n729), .EN(n218), .Y(a[2]) );
  TBUFX2 \myram/m12/ta/t1/b1  ( .A(n728), .EN(n218), .Y(a[1]) );
  TBUFX2 \myram/m12/ta/t0/b1  ( .A(n727), .EN(n218), .Y(a[0]) );
  TBUFX2 \myram/m11/tb/t31/b1  ( .A(n694), .EN(n257), .Y(b[31]) );
  TBUFX2 \myram/m11/tb/t30/b1  ( .A(n693), .EN(n257), .Y(b[30]) );
  TBUFX2 \myram/m11/tb/t29/b1  ( .A(n692), .EN(n257), .Y(b[29]) );
  TBUFX2 \myram/m11/tb/t28/b1  ( .A(n691), .EN(n257), .Y(b[28]) );
  TBUFX2 \myram/m11/tb/t27/b1  ( .A(n690), .EN(n257), .Y(b[27]) );
  TBUFX2 \myram/m11/tb/t26/b1  ( .A(n689), .EN(n257), .Y(b[26]) );
  TBUFX2 \myram/m11/tb/t25/b1  ( .A(n688), .EN(n257), .Y(b[25]) );
  TBUFX2 \myram/m11/tb/t24/b1  ( .A(n687), .EN(n257), .Y(b[24]) );
  TBUFX2 \myram/m11/tb/t23/b1  ( .A(n686), .EN(n257), .Y(b[23]) );
  TBUFX2 \myram/m11/tb/t22/b1  ( .A(n685), .EN(n257), .Y(b[22]) );
  TBUFX2 \myram/m11/tb/t21/b1  ( .A(n684), .EN(n257), .Y(b[21]) );
  TBUFX2 \myram/m11/tb/t20/b1  ( .A(n683), .EN(n257), .Y(b[20]) );
  TBUFX2 \myram/m11/tb/t19/b1  ( .A(n682), .EN(n257), .Y(b[19]) );
  TBUFX2 \myram/m11/tb/t18/b1  ( .A(n681), .EN(n257), .Y(b[18]) );
  TBUFX2 \myram/m11/tb/t17/b1  ( .A(n680), .EN(n257), .Y(b[17]) );
  TBUFX2 \myram/m11/tb/t16/b1  ( .A(n679), .EN(n257), .Y(b[16]) );
  TBUFX2 \myram/m11/tb/t15/b1  ( .A(n678), .EN(n257), .Y(b[15]) );
  TBUFX2 \myram/m11/tb/t14/b1  ( .A(n677), .EN(n257), .Y(b[14]) );
  TBUFX2 \myram/m11/tb/t13/b1  ( .A(n676), .EN(n257), .Y(b[13]) );
  TBUFX2 \myram/m11/tb/t12/b1  ( .A(n675), .EN(n256), .Y(b[12]) );
  TBUFX2 \myram/m11/tb/t11/b1  ( .A(n674), .EN(n256), .Y(b[11]) );
  TBUFX2 \myram/m11/tb/t10/b1  ( .A(n673), .EN(n256), .Y(b[10]) );
  TBUFX2 \myram/m11/tb/t9/b1  ( .A(n672), .EN(n256), .Y(b[9]) );
  TBUFX2 \myram/m11/tb/t8/b1  ( .A(n671), .EN(n256), .Y(b[8]) );
  TBUFX2 \myram/m11/tb/t7/b1  ( .A(n670), .EN(n256), .Y(b[7]) );
  TBUFX2 \myram/m11/tb/t6/b1  ( .A(n669), .EN(n256), .Y(b[6]) );
  TBUFX2 \myram/m11/tb/t5/b1  ( .A(n668), .EN(n256), .Y(b[5]) );
  INVX1 \myram/m11/tb/t4/U1  ( .A(\myram/m11/dout[4] ), .Y(n699) );
  TBUFX2 \myram/m11/tb/t4/b1  ( .A(n699), .EN(n256), .Y(b[4]) );
  INVX1 \myram/m11/tb/t3/U1  ( .A(\myram/m11/dout[3] ), .Y(n698) );
  TBUFX2 \myram/m11/tb/t3/b1  ( .A(n698), .EN(n256), .Y(b[3]) );
  INVX1 \myram/m11/tb/t2/U1  ( .A(\myram/m11/dout[2] ), .Y(n697) );
  TBUFX2 \myram/m11/tb/t2/b1  ( .A(n697), .EN(n256), .Y(b[2]) );
  INVX1 \myram/m11/tb/t1/U1  ( .A(\myram/m11/dout[1] ), .Y(n696) );
  TBUFX2 \myram/m11/tb/t1/b1  ( .A(n696), .EN(n256), .Y(b[1]) );
  INVX1 \myram/m11/tb/t0/U1  ( .A(\myram/m11/dout[0] ), .Y(n695) );
  TBUFX2 \myram/m11/tb/t0/b1  ( .A(n695), .EN(n256), .Y(b[0]) );
  INVX1 \myram/m11/ta/t31/U1  ( .A(\myram/m11/dout[31] ), .Y(n694) );
  TBUFX2 \myram/m11/ta/t31/b1  ( .A(n694), .EN(\myram/sel_a[11] ), .Y(a[31])
         );
  INVX1 \myram/m11/ta/t30/U1  ( .A(\myram/m11/dout[30] ), .Y(n693) );
  TBUFX2 \myram/m11/ta/t30/b1  ( .A(n693), .EN(\myram/sel_a[11] ), .Y(a[30])
         );
  INVX1 \myram/m11/ta/t29/U1  ( .A(\myram/m11/dout[29] ), .Y(n692) );
  TBUFX2 \myram/m11/ta/t29/b1  ( .A(n692), .EN(\myram/sel_a[11] ), .Y(a[29])
         );
  INVX1 \myram/m11/ta/t28/U1  ( .A(\myram/m11/dout[28] ), .Y(n691) );
  TBUFX2 \myram/m11/ta/t28/b1  ( .A(n691), .EN(\myram/sel_a[11] ), .Y(a[28])
         );
  INVX1 \myram/m11/ta/t27/U1  ( .A(\myram/m11/dout[27] ), .Y(n690) );
  TBUFX2 \myram/m11/ta/t27/b1  ( .A(n690), .EN(\myram/sel_a[11] ), .Y(a[27])
         );
  INVX1 \myram/m11/ta/t26/U1  ( .A(\myram/m11/dout[26] ), .Y(n689) );
  TBUFX2 \myram/m11/ta/t26/b1  ( .A(n689), .EN(\myram/sel_a[11] ), .Y(a[26])
         );
  INVX1 \myram/m11/ta/t25/U1  ( .A(\myram/m11/dout[25] ), .Y(n688) );
  TBUFX2 \myram/m11/ta/t25/b1  ( .A(n688), .EN(\myram/sel_a[11] ), .Y(a[25])
         );
  INVX1 \myram/m11/ta/t24/U1  ( .A(\myram/m11/dout[24] ), .Y(n687) );
  TBUFX2 \myram/m11/ta/t24/b1  ( .A(n687), .EN(\myram/sel_a[11] ), .Y(a[24])
         );
  INVX1 \myram/m11/ta/t23/U1  ( .A(\myram/m11/dout[23] ), .Y(n686) );
  TBUFX2 \myram/m11/ta/t23/b1  ( .A(n686), .EN(\myram/sel_a[11] ), .Y(a[23])
         );
  INVX1 \myram/m11/ta/t22/U1  ( .A(\myram/m11/dout[22] ), .Y(n685) );
  TBUFX2 \myram/m11/ta/t22/b1  ( .A(n685), .EN(\myram/sel_a[11] ), .Y(a[22])
         );
  INVX1 \myram/m11/ta/t21/U1  ( .A(\myram/m11/dout[21] ), .Y(n684) );
  TBUFX2 \myram/m11/ta/t21/b1  ( .A(n684), .EN(\myram/sel_a[11] ), .Y(a[21])
         );
  INVX1 \myram/m11/ta/t20/U1  ( .A(\myram/m11/dout[20] ), .Y(n683) );
  TBUFX2 \myram/m11/ta/t20/b1  ( .A(n683), .EN(\myram/sel_a[11] ), .Y(a[20])
         );
  INVX1 \myram/m11/ta/t19/U1  ( .A(\myram/m11/dout[19] ), .Y(n682) );
  TBUFX2 \myram/m11/ta/t19/b1  ( .A(n682), .EN(\myram/sel_a[11] ), .Y(a[19])
         );
  INVX1 \myram/m11/ta/t18/U1  ( .A(\myram/m11/dout[18] ), .Y(n681) );
  TBUFX2 \myram/m11/ta/t18/b1  ( .A(n681), .EN(\myram/sel_a[11] ), .Y(a[18])
         );
  INVX1 \myram/m11/ta/t17/U1  ( .A(\myram/m11/dout[17] ), .Y(n680) );
  TBUFX2 \myram/m11/ta/t17/b1  ( .A(n680), .EN(\myram/sel_a[11] ), .Y(a[17])
         );
  INVX1 \myram/m11/ta/t16/U1  ( .A(\myram/m11/dout[16] ), .Y(n679) );
  TBUFX2 \myram/m11/ta/t16/b1  ( .A(n679), .EN(\myram/sel_a[11] ), .Y(a[16])
         );
  INVX1 \myram/m11/ta/t15/U1  ( .A(\myram/m11/dout[15] ), .Y(n678) );
  TBUFX2 \myram/m11/ta/t15/b1  ( .A(n678), .EN(\myram/sel_a[11] ), .Y(a[15])
         );
  INVX1 \myram/m11/ta/t14/U1  ( .A(\myram/m11/dout[14] ), .Y(n677) );
  TBUFX2 \myram/m11/ta/t14/b1  ( .A(n677), .EN(\myram/sel_a[11] ), .Y(a[14])
         );
  INVX1 \myram/m11/ta/t13/U1  ( .A(\myram/m11/dout[13] ), .Y(n676) );
  TBUFX2 \myram/m11/ta/t13/b1  ( .A(n676), .EN(n220), .Y(a[13]) );
  INVX1 \myram/m11/ta/t12/U1  ( .A(\myram/m11/dout[12] ), .Y(n675) );
  TBUFX2 \myram/m11/ta/t12/b1  ( .A(n675), .EN(n220), .Y(a[12]) );
  INVX1 \myram/m11/ta/t11/U1  ( .A(\myram/m11/dout[11] ), .Y(n674) );
  TBUFX2 \myram/m11/ta/t11/b1  ( .A(n674), .EN(n220), .Y(a[11]) );
  INVX1 \myram/m11/ta/t10/U1  ( .A(\myram/m11/dout[10] ), .Y(n673) );
  TBUFX2 \myram/m11/ta/t10/b1  ( .A(n673), .EN(n220), .Y(a[10]) );
  INVX1 \myram/m11/ta/t9/U1  ( .A(\myram/m11/dout[9] ), .Y(n672) );
  TBUFX2 \myram/m11/ta/t9/b1  ( .A(n672), .EN(n220), .Y(a[9]) );
  INVX1 \myram/m11/ta/t8/U1  ( .A(\myram/m11/dout[8] ), .Y(n671) );
  TBUFX2 \myram/m11/ta/t8/b1  ( .A(n671), .EN(n220), .Y(a[8]) );
  INVX1 \myram/m11/ta/t7/U1  ( .A(\myram/m11/dout[7] ), .Y(n670) );
  TBUFX2 \myram/m11/ta/t7/b1  ( .A(n670), .EN(n220), .Y(a[7]) );
  INVX1 \myram/m11/ta/t6/U1  ( .A(\myram/m11/dout[6] ), .Y(n669) );
  TBUFX2 \myram/m11/ta/t6/b1  ( .A(n669), .EN(n220), .Y(a[6]) );
  INVX1 \myram/m11/ta/t5/U1  ( .A(\myram/m11/dout[5] ), .Y(n668) );
  TBUFX2 \myram/m11/ta/t5/b1  ( .A(n668), .EN(n220), .Y(a[5]) );
  TBUFX2 \myram/m11/ta/t4/b1  ( .A(n699), .EN(n220), .Y(a[4]) );
  TBUFX2 \myram/m11/ta/t3/b1  ( .A(n698), .EN(n220), .Y(a[3]) );
  TBUFX2 \myram/m11/ta/t2/b1  ( .A(n697), .EN(n220), .Y(a[2]) );
  TBUFX2 \myram/m11/ta/t1/b1  ( .A(n696), .EN(n220), .Y(a[1]) );
  TBUFX2 \myram/m11/ta/t0/b1  ( .A(n695), .EN(n220), .Y(a[0]) );
  TBUFX2 \myram/m10/tb/t31/b1  ( .A(n662), .EN(n260), .Y(b[31]) );
  TBUFX2 \myram/m10/tb/t30/b1  ( .A(n661), .EN(n260), .Y(b[30]) );
  TBUFX2 \myram/m10/tb/t29/b1  ( .A(n660), .EN(n260), .Y(b[29]) );
  TBUFX2 \myram/m10/tb/t28/b1  ( .A(n659), .EN(n260), .Y(b[28]) );
  TBUFX2 \myram/m10/tb/t27/b1  ( .A(n658), .EN(n260), .Y(b[27]) );
  TBUFX2 \myram/m10/tb/t26/b1  ( .A(n657), .EN(n260), .Y(b[26]) );
  TBUFX2 \myram/m10/tb/t25/b1  ( .A(n656), .EN(n260), .Y(b[25]) );
  TBUFX2 \myram/m10/tb/t24/b1  ( .A(n655), .EN(n260), .Y(b[24]) );
  TBUFX2 \myram/m10/tb/t23/b1  ( .A(n654), .EN(n260), .Y(b[23]) );
  TBUFX2 \myram/m10/tb/t22/b1  ( .A(n653), .EN(n260), .Y(b[22]) );
  TBUFX2 \myram/m10/tb/t21/b1  ( .A(n652), .EN(n260), .Y(b[21]) );
  TBUFX2 \myram/m10/tb/t20/b1  ( .A(n651), .EN(n260), .Y(b[20]) );
  TBUFX2 \myram/m10/tb/t19/b1  ( .A(n650), .EN(n260), .Y(b[19]) );
  TBUFX2 \myram/m10/tb/t18/b1  ( .A(n649), .EN(n260), .Y(b[18]) );
  TBUFX2 \myram/m10/tb/t17/b1  ( .A(n648), .EN(n260), .Y(b[17]) );
  TBUFX2 \myram/m10/tb/t16/b1  ( .A(n647), .EN(n260), .Y(b[16]) );
  TBUFX2 \myram/m10/tb/t15/b1  ( .A(n646), .EN(n260), .Y(b[15]) );
  TBUFX2 \myram/m10/tb/t14/b1  ( .A(n645), .EN(n260), .Y(b[14]) );
  TBUFX2 \myram/m10/tb/t13/b1  ( .A(n644), .EN(n260), .Y(b[13]) );
  TBUFX2 \myram/m10/tb/t12/b1  ( .A(n643), .EN(n259), .Y(b[12]) );
  TBUFX2 \myram/m10/tb/t11/b1  ( .A(n642), .EN(n259), .Y(b[11]) );
  TBUFX2 \myram/m10/tb/t10/b1  ( .A(n641), .EN(n259), .Y(b[10]) );
  TBUFX2 \myram/m10/tb/t9/b1  ( .A(n640), .EN(n259), .Y(b[9]) );
  TBUFX2 \myram/m10/tb/t8/b1  ( .A(n639), .EN(n259), .Y(b[8]) );
  TBUFX2 \myram/m10/tb/t7/b1  ( .A(n638), .EN(n259), .Y(b[7]) );
  TBUFX2 \myram/m10/tb/t6/b1  ( .A(n637), .EN(n259), .Y(b[6]) );
  TBUFX2 \myram/m10/tb/t5/b1  ( .A(n636), .EN(n259), .Y(b[5]) );
  INVX1 \myram/m10/tb/t4/U1  ( .A(\myram/m10/dout[4] ), .Y(n667) );
  TBUFX2 \myram/m10/tb/t4/b1  ( .A(n667), .EN(n259), .Y(b[4]) );
  INVX1 \myram/m10/tb/t3/U1  ( .A(\myram/m10/dout[3] ), .Y(n666) );
  TBUFX2 \myram/m10/tb/t3/b1  ( .A(n666), .EN(n259), .Y(b[3]) );
  INVX1 \myram/m10/tb/t2/U1  ( .A(\myram/m10/dout[2] ), .Y(n665) );
  TBUFX2 \myram/m10/tb/t2/b1  ( .A(n665), .EN(n259), .Y(b[2]) );
  INVX1 \myram/m10/tb/t1/U1  ( .A(\myram/m10/dout[1] ), .Y(n664) );
  TBUFX2 \myram/m10/tb/t1/b1  ( .A(n664), .EN(n259), .Y(b[1]) );
  INVX1 \myram/m10/tb/t0/U1  ( .A(\myram/m10/dout[0] ), .Y(n663) );
  TBUFX2 \myram/m10/tb/t0/b1  ( .A(n663), .EN(n259), .Y(b[0]) );
  INVX1 \myram/m10/ta/t31/U1  ( .A(\myram/m10/dout[31] ), .Y(n662) );
  TBUFX2 \myram/m10/ta/t31/b1  ( .A(n662), .EN(\myram/sel_a[10] ), .Y(a[31])
         );
  INVX1 \myram/m10/ta/t30/U1  ( .A(\myram/m10/dout[30] ), .Y(n661) );
  TBUFX2 \myram/m10/ta/t30/b1  ( .A(n661), .EN(\myram/sel_a[10] ), .Y(a[30])
         );
  INVX1 \myram/m10/ta/t29/U1  ( .A(\myram/m10/dout[29] ), .Y(n660) );
  TBUFX2 \myram/m10/ta/t29/b1  ( .A(n660), .EN(\myram/sel_a[10] ), .Y(a[29])
         );
  INVX1 \myram/m10/ta/t28/U1  ( .A(\myram/m10/dout[28] ), .Y(n659) );
  TBUFX2 \myram/m10/ta/t28/b1  ( .A(n659), .EN(\myram/sel_a[10] ), .Y(a[28])
         );
  INVX1 \myram/m10/ta/t27/U1  ( .A(\myram/m10/dout[27] ), .Y(n658) );
  TBUFX2 \myram/m10/ta/t27/b1  ( .A(n658), .EN(\myram/sel_a[10] ), .Y(a[27])
         );
  INVX1 \myram/m10/ta/t26/U1  ( .A(\myram/m10/dout[26] ), .Y(n657) );
  TBUFX2 \myram/m10/ta/t26/b1  ( .A(n657), .EN(\myram/sel_a[10] ), .Y(a[26])
         );
  INVX1 \myram/m10/ta/t25/U1  ( .A(\myram/m10/dout[25] ), .Y(n656) );
  TBUFX2 \myram/m10/ta/t25/b1  ( .A(n656), .EN(\myram/sel_a[10] ), .Y(a[25])
         );
  INVX1 \myram/m10/ta/t24/U1  ( .A(\myram/m10/dout[24] ), .Y(n655) );
  TBUFX2 \myram/m10/ta/t24/b1  ( .A(n655), .EN(\myram/sel_a[10] ), .Y(a[24])
         );
  INVX1 \myram/m10/ta/t23/U1  ( .A(\myram/m10/dout[23] ), .Y(n654) );
  TBUFX2 \myram/m10/ta/t23/b1  ( .A(n654), .EN(\myram/sel_a[10] ), .Y(a[23])
         );
  INVX1 \myram/m10/ta/t22/U1  ( .A(\myram/m10/dout[22] ), .Y(n653) );
  TBUFX2 \myram/m10/ta/t22/b1  ( .A(n653), .EN(\myram/sel_a[10] ), .Y(a[22])
         );
  INVX1 \myram/m10/ta/t21/U1  ( .A(\myram/m10/dout[21] ), .Y(n652) );
  TBUFX2 \myram/m10/ta/t21/b1  ( .A(n652), .EN(\myram/sel_a[10] ), .Y(a[21])
         );
  INVX1 \myram/m10/ta/t20/U1  ( .A(\myram/m10/dout[20] ), .Y(n651) );
  TBUFX2 \myram/m10/ta/t20/b1  ( .A(n651), .EN(\myram/sel_a[10] ), .Y(a[20])
         );
  INVX1 \myram/m10/ta/t19/U1  ( .A(\myram/m10/dout[19] ), .Y(n650) );
  TBUFX2 \myram/m10/ta/t19/b1  ( .A(n650), .EN(\myram/sel_a[10] ), .Y(a[19])
         );
  INVX1 \myram/m10/ta/t18/U1  ( .A(\myram/m10/dout[18] ), .Y(n649) );
  TBUFX2 \myram/m10/ta/t18/b1  ( .A(n649), .EN(\myram/sel_a[10] ), .Y(a[18])
         );
  INVX1 \myram/m10/ta/t17/U1  ( .A(\myram/m10/dout[17] ), .Y(n648) );
  TBUFX2 \myram/m10/ta/t17/b1  ( .A(n648), .EN(\myram/sel_a[10] ), .Y(a[17])
         );
  INVX1 \myram/m10/ta/t16/U1  ( .A(\myram/m10/dout[16] ), .Y(n647) );
  TBUFX2 \myram/m10/ta/t16/b1  ( .A(n647), .EN(\myram/sel_a[10] ), .Y(a[16])
         );
  INVX1 \myram/m10/ta/t15/U1  ( .A(\myram/m10/dout[15] ), .Y(n646) );
  TBUFX2 \myram/m10/ta/t15/b1  ( .A(n646), .EN(\myram/sel_a[10] ), .Y(a[15])
         );
  INVX1 \myram/m10/ta/t14/U1  ( .A(\myram/m10/dout[14] ), .Y(n645) );
  TBUFX2 \myram/m10/ta/t14/b1  ( .A(n645), .EN(\myram/sel_a[10] ), .Y(a[14])
         );
  INVX1 \myram/m10/ta/t13/U1  ( .A(\myram/m10/dout[13] ), .Y(n644) );
  TBUFX2 \myram/m10/ta/t13/b1  ( .A(n644), .EN(n222), .Y(a[13]) );
  INVX1 \myram/m10/ta/t12/U1  ( .A(\myram/m10/dout[12] ), .Y(n643) );
  TBUFX2 \myram/m10/ta/t12/b1  ( .A(n643), .EN(n222), .Y(a[12]) );
  INVX1 \myram/m10/ta/t11/U1  ( .A(\myram/m10/dout[11] ), .Y(n642) );
  TBUFX2 \myram/m10/ta/t11/b1  ( .A(n642), .EN(n222), .Y(a[11]) );
  INVX1 \myram/m10/ta/t10/U1  ( .A(\myram/m10/dout[10] ), .Y(n641) );
  TBUFX2 \myram/m10/ta/t10/b1  ( .A(n641), .EN(n222), .Y(a[10]) );
  INVX1 \myram/m10/ta/t9/U1  ( .A(\myram/m10/dout[9] ), .Y(n640) );
  TBUFX2 \myram/m10/ta/t9/b1  ( .A(n640), .EN(n222), .Y(a[9]) );
  INVX1 \myram/m10/ta/t8/U1  ( .A(\myram/m10/dout[8] ), .Y(n639) );
  TBUFX2 \myram/m10/ta/t8/b1  ( .A(n639), .EN(n222), .Y(a[8]) );
  INVX1 \myram/m10/ta/t7/U1  ( .A(\myram/m10/dout[7] ), .Y(n638) );
  TBUFX2 \myram/m10/ta/t7/b1  ( .A(n638), .EN(n222), .Y(a[7]) );
  INVX1 \myram/m10/ta/t6/U1  ( .A(\myram/m10/dout[6] ), .Y(n637) );
  TBUFX2 \myram/m10/ta/t6/b1  ( .A(n637), .EN(n222), .Y(a[6]) );
  INVX1 \myram/m10/ta/t5/U1  ( .A(\myram/m10/dout[5] ), .Y(n636) );
  TBUFX2 \myram/m10/ta/t5/b1  ( .A(n636), .EN(n222), .Y(a[5]) );
  TBUFX2 \myram/m10/ta/t4/b1  ( .A(n667), .EN(n222), .Y(a[4]) );
  TBUFX2 \myram/m10/ta/t3/b1  ( .A(n666), .EN(n222), .Y(a[3]) );
  TBUFX2 \myram/m10/ta/t2/b1  ( .A(n665), .EN(n222), .Y(a[2]) );
  TBUFX2 \myram/m10/ta/t1/b1  ( .A(n664), .EN(n222), .Y(a[1]) );
  TBUFX2 \myram/m10/ta/t0/b1  ( .A(n663), .EN(n222), .Y(a[0]) );
  TBUFX2 \myram/m9/tb/t31/b1  ( .A(n630), .EN(n263), .Y(b[31]) );
  TBUFX2 \myram/m9/tb/t30/b1  ( .A(n629), .EN(n263), .Y(b[30]) );
  TBUFX2 \myram/m9/tb/t29/b1  ( .A(n628), .EN(n263), .Y(b[29]) );
  TBUFX2 \myram/m9/tb/t28/b1  ( .A(n627), .EN(n263), .Y(b[28]) );
  TBUFX2 \myram/m9/tb/t27/b1  ( .A(n626), .EN(n263), .Y(b[27]) );
  TBUFX2 \myram/m9/tb/t26/b1  ( .A(n625), .EN(n263), .Y(b[26]) );
  TBUFX2 \myram/m9/tb/t25/b1  ( .A(n624), .EN(n263), .Y(b[25]) );
  TBUFX2 \myram/m9/tb/t24/b1  ( .A(n623), .EN(n263), .Y(b[24]) );
  TBUFX2 \myram/m9/tb/t23/b1  ( .A(n622), .EN(n263), .Y(b[23]) );
  TBUFX2 \myram/m9/tb/t22/b1  ( .A(n621), .EN(n263), .Y(b[22]) );
  TBUFX2 \myram/m9/tb/t21/b1  ( .A(n620), .EN(n263), .Y(b[21]) );
  TBUFX2 \myram/m9/tb/t20/b1  ( .A(n619), .EN(n263), .Y(b[20]) );
  TBUFX2 \myram/m9/tb/t19/b1  ( .A(n618), .EN(n263), .Y(b[19]) );
  TBUFX2 \myram/m9/tb/t18/b1  ( .A(n617), .EN(n263), .Y(b[18]) );
  TBUFX2 \myram/m9/tb/t17/b1  ( .A(n616), .EN(n263), .Y(b[17]) );
  TBUFX2 \myram/m9/tb/t16/b1  ( .A(n615), .EN(n263), .Y(b[16]) );
  TBUFX2 \myram/m9/tb/t15/b1  ( .A(n614), .EN(n263), .Y(b[15]) );
  TBUFX2 \myram/m9/tb/t14/b1  ( .A(n613), .EN(n263), .Y(b[14]) );
  TBUFX2 \myram/m9/tb/t13/b1  ( .A(n612), .EN(n263), .Y(b[13]) );
  TBUFX2 \myram/m9/tb/t12/b1  ( .A(n611), .EN(n262), .Y(b[12]) );
  TBUFX2 \myram/m9/tb/t11/b1  ( .A(n610), .EN(n262), .Y(b[11]) );
  TBUFX2 \myram/m9/tb/t10/b1  ( .A(n609), .EN(n262), .Y(b[10]) );
  TBUFX2 \myram/m9/tb/t9/b1  ( .A(n608), .EN(n262), .Y(b[9]) );
  TBUFX2 \myram/m9/tb/t8/b1  ( .A(n607), .EN(n262), .Y(b[8]) );
  TBUFX2 \myram/m9/tb/t7/b1  ( .A(n606), .EN(n262), .Y(b[7]) );
  TBUFX2 \myram/m9/tb/t6/b1  ( .A(n605), .EN(n262), .Y(b[6]) );
  TBUFX2 \myram/m9/tb/t5/b1  ( .A(n604), .EN(n262), .Y(b[5]) );
  INVX1 \myram/m9/tb/t4/U1  ( .A(\myram/m9/dout[4] ), .Y(n635) );
  TBUFX2 \myram/m9/tb/t4/b1  ( .A(n635), .EN(n262), .Y(b[4]) );
  INVX1 \myram/m9/tb/t3/U1  ( .A(\myram/m9/dout[3] ), .Y(n634) );
  TBUFX2 \myram/m9/tb/t3/b1  ( .A(n634), .EN(n262), .Y(b[3]) );
  INVX1 \myram/m9/tb/t2/U1  ( .A(\myram/m9/dout[2] ), .Y(n633) );
  TBUFX2 \myram/m9/tb/t2/b1  ( .A(n633), .EN(n262), .Y(b[2]) );
  INVX1 \myram/m9/tb/t1/U1  ( .A(\myram/m9/dout[1] ), .Y(n632) );
  TBUFX2 \myram/m9/tb/t1/b1  ( .A(n632), .EN(n262), .Y(b[1]) );
  INVX1 \myram/m9/tb/t0/U1  ( .A(\myram/m9/dout[0] ), .Y(n631) );
  TBUFX2 \myram/m9/tb/t0/b1  ( .A(n631), .EN(n262), .Y(b[0]) );
  INVX1 \myram/m9/ta/t31/U1  ( .A(\myram/m9/dout[31] ), .Y(n630) );
  TBUFX2 \myram/m9/ta/t31/b1  ( .A(n630), .EN(\myram/sel_a[9] ), .Y(a[31]) );
  INVX1 \myram/m9/ta/t30/U1  ( .A(\myram/m9/dout[30] ), .Y(n629) );
  TBUFX2 \myram/m9/ta/t30/b1  ( .A(n629), .EN(\myram/sel_a[9] ), .Y(a[30]) );
  INVX1 \myram/m9/ta/t29/U1  ( .A(\myram/m9/dout[29] ), .Y(n628) );
  TBUFX2 \myram/m9/ta/t29/b1  ( .A(n628), .EN(\myram/sel_a[9] ), .Y(a[29]) );
  INVX1 \myram/m9/ta/t28/U1  ( .A(\myram/m9/dout[28] ), .Y(n627) );
  TBUFX2 \myram/m9/ta/t28/b1  ( .A(n627), .EN(\myram/sel_a[9] ), .Y(a[28]) );
  INVX1 \myram/m9/ta/t27/U1  ( .A(\myram/m9/dout[27] ), .Y(n626) );
  TBUFX2 \myram/m9/ta/t27/b1  ( .A(n626), .EN(\myram/sel_a[9] ), .Y(a[27]) );
  INVX1 \myram/m9/ta/t26/U1  ( .A(\myram/m9/dout[26] ), .Y(n625) );
  TBUFX2 \myram/m9/ta/t26/b1  ( .A(n625), .EN(\myram/sel_a[9] ), .Y(a[26]) );
  INVX1 \myram/m9/ta/t25/U1  ( .A(\myram/m9/dout[25] ), .Y(n624) );
  TBUFX2 \myram/m9/ta/t25/b1  ( .A(n624), .EN(\myram/sel_a[9] ), .Y(a[25]) );
  INVX1 \myram/m9/ta/t24/U1  ( .A(\myram/m9/dout[24] ), .Y(n623) );
  TBUFX2 \myram/m9/ta/t24/b1  ( .A(n623), .EN(\myram/sel_a[9] ), .Y(a[24]) );
  INVX1 \myram/m9/ta/t23/U1  ( .A(\myram/m9/dout[23] ), .Y(n622) );
  TBUFX2 \myram/m9/ta/t23/b1  ( .A(n622), .EN(\myram/sel_a[9] ), .Y(a[23]) );
  INVX1 \myram/m9/ta/t22/U1  ( .A(\myram/m9/dout[22] ), .Y(n621) );
  TBUFX2 \myram/m9/ta/t22/b1  ( .A(n621), .EN(\myram/sel_a[9] ), .Y(a[22]) );
  INVX1 \myram/m9/ta/t21/U1  ( .A(\myram/m9/dout[21] ), .Y(n620) );
  TBUFX2 \myram/m9/ta/t21/b1  ( .A(n620), .EN(\myram/sel_a[9] ), .Y(a[21]) );
  INVX1 \myram/m9/ta/t20/U1  ( .A(\myram/m9/dout[20] ), .Y(n619) );
  TBUFX2 \myram/m9/ta/t20/b1  ( .A(n619), .EN(\myram/sel_a[9] ), .Y(a[20]) );
  INVX1 \myram/m9/ta/t19/U1  ( .A(\myram/m9/dout[19] ), .Y(n618) );
  TBUFX2 \myram/m9/ta/t19/b1  ( .A(n618), .EN(\myram/sel_a[9] ), .Y(a[19]) );
  INVX1 \myram/m9/ta/t18/U1  ( .A(\myram/m9/dout[18] ), .Y(n617) );
  TBUFX2 \myram/m9/ta/t18/b1  ( .A(n617), .EN(\myram/sel_a[9] ), .Y(a[18]) );
  INVX1 \myram/m9/ta/t17/U1  ( .A(\myram/m9/dout[17] ), .Y(n616) );
  TBUFX2 \myram/m9/ta/t17/b1  ( .A(n616), .EN(\myram/sel_a[9] ), .Y(a[17]) );
  INVX1 \myram/m9/ta/t16/U1  ( .A(\myram/m9/dout[16] ), .Y(n615) );
  TBUFX2 \myram/m9/ta/t16/b1  ( .A(n615), .EN(\myram/sel_a[9] ), .Y(a[16]) );
  INVX1 \myram/m9/ta/t15/U1  ( .A(\myram/m9/dout[15] ), .Y(n614) );
  TBUFX2 \myram/m9/ta/t15/b1  ( .A(n614), .EN(\myram/sel_a[9] ), .Y(a[15]) );
  INVX1 \myram/m9/ta/t14/U1  ( .A(\myram/m9/dout[14] ), .Y(n613) );
  TBUFX2 \myram/m9/ta/t14/b1  ( .A(n613), .EN(\myram/sel_a[9] ), .Y(a[14]) );
  INVX1 \myram/m9/ta/t13/U1  ( .A(\myram/m9/dout[13] ), .Y(n612) );
  TBUFX2 \myram/m9/ta/t13/b1  ( .A(n612), .EN(n224), .Y(a[13]) );
  INVX1 \myram/m9/ta/t12/U1  ( .A(\myram/m9/dout[12] ), .Y(n611) );
  TBUFX2 \myram/m9/ta/t12/b1  ( .A(n611), .EN(n224), .Y(a[12]) );
  INVX1 \myram/m9/ta/t11/U1  ( .A(\myram/m9/dout[11] ), .Y(n610) );
  TBUFX2 \myram/m9/ta/t11/b1  ( .A(n610), .EN(n224), .Y(a[11]) );
  INVX1 \myram/m9/ta/t10/U1  ( .A(\myram/m9/dout[10] ), .Y(n609) );
  TBUFX2 \myram/m9/ta/t10/b1  ( .A(n609), .EN(n224), .Y(a[10]) );
  INVX1 \myram/m9/ta/t9/U1  ( .A(\myram/m9/dout[9] ), .Y(n608) );
  TBUFX2 \myram/m9/ta/t9/b1  ( .A(n608), .EN(n224), .Y(a[9]) );
  INVX1 \myram/m9/ta/t8/U1  ( .A(\myram/m9/dout[8] ), .Y(n607) );
  TBUFX2 \myram/m9/ta/t8/b1  ( .A(n607), .EN(n224), .Y(a[8]) );
  INVX1 \myram/m9/ta/t7/U1  ( .A(\myram/m9/dout[7] ), .Y(n606) );
  TBUFX2 \myram/m9/ta/t7/b1  ( .A(n606), .EN(n224), .Y(a[7]) );
  INVX1 \myram/m9/ta/t6/U1  ( .A(\myram/m9/dout[6] ), .Y(n605) );
  TBUFX2 \myram/m9/ta/t6/b1  ( .A(n605), .EN(n224), .Y(a[6]) );
  INVX1 \myram/m9/ta/t5/U1  ( .A(\myram/m9/dout[5] ), .Y(n604) );
  TBUFX2 \myram/m9/ta/t5/b1  ( .A(n604), .EN(n224), .Y(a[5]) );
  TBUFX2 \myram/m9/ta/t4/b1  ( .A(n635), .EN(n224), .Y(a[4]) );
  TBUFX2 \myram/m9/ta/t3/b1  ( .A(n634), .EN(n224), .Y(a[3]) );
  TBUFX2 \myram/m9/ta/t2/b1  ( .A(n633), .EN(n224), .Y(a[2]) );
  TBUFX2 \myram/m9/ta/t1/b1  ( .A(n632), .EN(n224), .Y(a[1]) );
  TBUFX2 \myram/m9/ta/t0/b1  ( .A(n631), .EN(n224), .Y(a[0]) );
  TBUFX2 \myram/m8/tb/t31/b1  ( .A(n598), .EN(n266), .Y(b[31]) );
  TBUFX2 \myram/m8/tb/t30/b1  ( .A(n597), .EN(n266), .Y(b[30]) );
  TBUFX2 \myram/m8/tb/t29/b1  ( .A(n596), .EN(n266), .Y(b[29]) );
  TBUFX2 \myram/m8/tb/t28/b1  ( .A(n595), .EN(n266), .Y(b[28]) );
  TBUFX2 \myram/m8/tb/t27/b1  ( .A(n594), .EN(n266), .Y(b[27]) );
  TBUFX2 \myram/m8/tb/t26/b1  ( .A(n593), .EN(n266), .Y(b[26]) );
  TBUFX2 \myram/m8/tb/t25/b1  ( .A(n592), .EN(n266), .Y(b[25]) );
  TBUFX2 \myram/m8/tb/t24/b1  ( .A(n591), .EN(n266), .Y(b[24]) );
  TBUFX2 \myram/m8/tb/t23/b1  ( .A(n590), .EN(n266), .Y(b[23]) );
  TBUFX2 \myram/m8/tb/t22/b1  ( .A(n589), .EN(n266), .Y(b[22]) );
  TBUFX2 \myram/m8/tb/t21/b1  ( .A(n588), .EN(n266), .Y(b[21]) );
  TBUFX2 \myram/m8/tb/t20/b1  ( .A(n587), .EN(n266), .Y(b[20]) );
  TBUFX2 \myram/m8/tb/t19/b1  ( .A(n586), .EN(n266), .Y(b[19]) );
  TBUFX2 \myram/m8/tb/t18/b1  ( .A(n585), .EN(n266), .Y(b[18]) );
  TBUFX2 \myram/m8/tb/t17/b1  ( .A(n584), .EN(n266), .Y(b[17]) );
  TBUFX2 \myram/m8/tb/t16/b1  ( .A(n583), .EN(n266), .Y(b[16]) );
  TBUFX2 \myram/m8/tb/t15/b1  ( .A(n582), .EN(n266), .Y(b[15]) );
  TBUFX2 \myram/m8/tb/t14/b1  ( .A(n581), .EN(n266), .Y(b[14]) );
  TBUFX2 \myram/m8/tb/t13/b1  ( .A(n580), .EN(n266), .Y(b[13]) );
  TBUFX2 \myram/m8/tb/t12/b1  ( .A(n579), .EN(n265), .Y(b[12]) );
  TBUFX2 \myram/m8/tb/t11/b1  ( .A(n578), .EN(n265), .Y(b[11]) );
  TBUFX2 \myram/m8/tb/t10/b1  ( .A(n577), .EN(n265), .Y(b[10]) );
  TBUFX2 \myram/m8/tb/t9/b1  ( .A(n576), .EN(n265), .Y(b[9]) );
  TBUFX2 \myram/m8/tb/t8/b1  ( .A(n575), .EN(n265), .Y(b[8]) );
  TBUFX2 \myram/m8/tb/t7/b1  ( .A(n574), .EN(n265), .Y(b[7]) );
  TBUFX2 \myram/m8/tb/t6/b1  ( .A(n573), .EN(n265), .Y(b[6]) );
  TBUFX2 \myram/m8/tb/t5/b1  ( .A(n572), .EN(n265), .Y(b[5]) );
  INVX1 \myram/m8/tb/t4/U1  ( .A(\myram/m8/dout[4] ), .Y(n603) );
  TBUFX2 \myram/m8/tb/t4/b1  ( .A(n603), .EN(n265), .Y(b[4]) );
  INVX1 \myram/m8/tb/t3/U1  ( .A(\myram/m8/dout[3] ), .Y(n602) );
  TBUFX2 \myram/m8/tb/t3/b1  ( .A(n602), .EN(n265), .Y(b[3]) );
  INVX1 \myram/m8/tb/t2/U1  ( .A(\myram/m8/dout[2] ), .Y(n601) );
  TBUFX2 \myram/m8/tb/t2/b1  ( .A(n601), .EN(n265), .Y(b[2]) );
  INVX1 \myram/m8/tb/t1/U1  ( .A(\myram/m8/dout[1] ), .Y(n600) );
  TBUFX2 \myram/m8/tb/t1/b1  ( .A(n600), .EN(n265), .Y(b[1]) );
  INVX1 \myram/m8/tb/t0/U1  ( .A(\myram/m8/dout[0] ), .Y(n599) );
  TBUFX2 \myram/m8/tb/t0/b1  ( .A(n599), .EN(n265), .Y(b[0]) );
  INVX1 \myram/m8/ta/t31/U1  ( .A(\myram/m8/dout[31] ), .Y(n598) );
  TBUFX2 \myram/m8/ta/t31/b1  ( .A(n598), .EN(\myram/sel_a[8] ), .Y(a[31]) );
  INVX1 \myram/m8/ta/t30/U1  ( .A(\myram/m8/dout[30] ), .Y(n597) );
  TBUFX2 \myram/m8/ta/t30/b1  ( .A(n597), .EN(\myram/sel_a[8] ), .Y(a[30]) );
  INVX1 \myram/m8/ta/t29/U1  ( .A(\myram/m8/dout[29] ), .Y(n596) );
  TBUFX2 \myram/m8/ta/t29/b1  ( .A(n596), .EN(\myram/sel_a[8] ), .Y(a[29]) );
  INVX1 \myram/m8/ta/t28/U1  ( .A(\myram/m8/dout[28] ), .Y(n595) );
  TBUFX2 \myram/m8/ta/t28/b1  ( .A(n595), .EN(\myram/sel_a[8] ), .Y(a[28]) );
  INVX1 \myram/m8/ta/t27/U1  ( .A(\myram/m8/dout[27] ), .Y(n594) );
  TBUFX2 \myram/m8/ta/t27/b1  ( .A(n594), .EN(\myram/sel_a[8] ), .Y(a[27]) );
  INVX1 \myram/m8/ta/t26/U1  ( .A(\myram/m8/dout[26] ), .Y(n593) );
  TBUFX2 \myram/m8/ta/t26/b1  ( .A(n593), .EN(\myram/sel_a[8] ), .Y(a[26]) );
  INVX1 \myram/m8/ta/t25/U1  ( .A(\myram/m8/dout[25] ), .Y(n592) );
  TBUFX2 \myram/m8/ta/t25/b1  ( .A(n592), .EN(\myram/sel_a[8] ), .Y(a[25]) );
  INVX1 \myram/m8/ta/t24/U1  ( .A(\myram/m8/dout[24] ), .Y(n591) );
  TBUFX2 \myram/m8/ta/t24/b1  ( .A(n591), .EN(\myram/sel_a[8] ), .Y(a[24]) );
  INVX1 \myram/m8/ta/t23/U1  ( .A(\myram/m8/dout[23] ), .Y(n590) );
  TBUFX2 \myram/m8/ta/t23/b1  ( .A(n590), .EN(\myram/sel_a[8] ), .Y(a[23]) );
  INVX1 \myram/m8/ta/t22/U1  ( .A(\myram/m8/dout[22] ), .Y(n589) );
  TBUFX2 \myram/m8/ta/t22/b1  ( .A(n589), .EN(\myram/sel_a[8] ), .Y(a[22]) );
  INVX1 \myram/m8/ta/t21/U1  ( .A(\myram/m8/dout[21] ), .Y(n588) );
  TBUFX2 \myram/m8/ta/t21/b1  ( .A(n588), .EN(\myram/sel_a[8] ), .Y(a[21]) );
  INVX1 \myram/m8/ta/t20/U1  ( .A(\myram/m8/dout[20] ), .Y(n587) );
  TBUFX2 \myram/m8/ta/t20/b1  ( .A(n587), .EN(\myram/sel_a[8] ), .Y(a[20]) );
  INVX1 \myram/m8/ta/t19/U1  ( .A(\myram/m8/dout[19] ), .Y(n586) );
  TBUFX2 \myram/m8/ta/t19/b1  ( .A(n586), .EN(\myram/sel_a[8] ), .Y(a[19]) );
  INVX1 \myram/m8/ta/t18/U1  ( .A(\myram/m8/dout[18] ), .Y(n585) );
  TBUFX2 \myram/m8/ta/t18/b1  ( .A(n585), .EN(\myram/sel_a[8] ), .Y(a[18]) );
  INVX1 \myram/m8/ta/t17/U1  ( .A(\myram/m8/dout[17] ), .Y(n584) );
  TBUFX2 \myram/m8/ta/t17/b1  ( .A(n584), .EN(\myram/sel_a[8] ), .Y(a[17]) );
  INVX1 \myram/m8/ta/t16/U1  ( .A(\myram/m8/dout[16] ), .Y(n583) );
  TBUFX2 \myram/m8/ta/t16/b1  ( .A(n583), .EN(\myram/sel_a[8] ), .Y(a[16]) );
  INVX1 \myram/m8/ta/t15/U1  ( .A(\myram/m8/dout[15] ), .Y(n582) );
  TBUFX2 \myram/m8/ta/t15/b1  ( .A(n582), .EN(\myram/sel_a[8] ), .Y(a[15]) );
  INVX1 \myram/m8/ta/t14/U1  ( .A(\myram/m8/dout[14] ), .Y(n581) );
  TBUFX2 \myram/m8/ta/t14/b1  ( .A(n581), .EN(\myram/sel_a[8] ), .Y(a[14]) );
  INVX1 \myram/m8/ta/t13/U1  ( .A(\myram/m8/dout[13] ), .Y(n580) );
  TBUFX2 \myram/m8/ta/t13/b1  ( .A(n580), .EN(n226), .Y(a[13]) );
  INVX1 \myram/m8/ta/t12/U1  ( .A(\myram/m8/dout[12] ), .Y(n579) );
  TBUFX2 \myram/m8/ta/t12/b1  ( .A(n579), .EN(n226), .Y(a[12]) );
  INVX1 \myram/m8/ta/t11/U1  ( .A(\myram/m8/dout[11] ), .Y(n578) );
  TBUFX2 \myram/m8/ta/t11/b1  ( .A(n578), .EN(n226), .Y(a[11]) );
  INVX1 \myram/m8/ta/t10/U1  ( .A(\myram/m8/dout[10] ), .Y(n577) );
  TBUFX2 \myram/m8/ta/t10/b1  ( .A(n577), .EN(n226), .Y(a[10]) );
  INVX1 \myram/m8/ta/t9/U1  ( .A(\myram/m8/dout[9] ), .Y(n576) );
  TBUFX2 \myram/m8/ta/t9/b1  ( .A(n576), .EN(n226), .Y(a[9]) );
  INVX1 \myram/m8/ta/t8/U1  ( .A(\myram/m8/dout[8] ), .Y(n575) );
  TBUFX2 \myram/m8/ta/t8/b1  ( .A(n575), .EN(n226), .Y(a[8]) );
  INVX1 \myram/m8/ta/t7/U1  ( .A(\myram/m8/dout[7] ), .Y(n574) );
  TBUFX2 \myram/m8/ta/t7/b1  ( .A(n574), .EN(n226), .Y(a[7]) );
  INVX1 \myram/m8/ta/t6/U1  ( .A(\myram/m8/dout[6] ), .Y(n573) );
  TBUFX2 \myram/m8/ta/t6/b1  ( .A(n573), .EN(n226), .Y(a[6]) );
  INVX1 \myram/m8/ta/t5/U1  ( .A(\myram/m8/dout[5] ), .Y(n572) );
  TBUFX2 \myram/m8/ta/t5/b1  ( .A(n572), .EN(n226), .Y(a[5]) );
  TBUFX2 \myram/m8/ta/t4/b1  ( .A(n603), .EN(n226), .Y(a[4]) );
  TBUFX2 \myram/m8/ta/t3/b1  ( .A(n602), .EN(n226), .Y(a[3]) );
  TBUFX2 \myram/m8/ta/t2/b1  ( .A(n601), .EN(n226), .Y(a[2]) );
  TBUFX2 \myram/m8/ta/t1/b1  ( .A(n600), .EN(n226), .Y(a[1]) );
  TBUFX2 \myram/m8/ta/t0/b1  ( .A(n599), .EN(n226), .Y(a[0]) );
  TBUFX2 \myram/m7/tb/t31/b1  ( .A(n566), .EN(n269), .Y(b[31]) );
  TBUFX2 \myram/m7/tb/t30/b1  ( .A(n565), .EN(n269), .Y(b[30]) );
  TBUFX2 \myram/m7/tb/t29/b1  ( .A(n564), .EN(n269), .Y(b[29]) );
  TBUFX2 \myram/m7/tb/t28/b1  ( .A(n563), .EN(n269), .Y(b[28]) );
  TBUFX2 \myram/m7/tb/t27/b1  ( .A(n562), .EN(n269), .Y(b[27]) );
  TBUFX2 \myram/m7/tb/t26/b1  ( .A(n561), .EN(n269), .Y(b[26]) );
  TBUFX2 \myram/m7/tb/t25/b1  ( .A(n560), .EN(n269), .Y(b[25]) );
  TBUFX2 \myram/m7/tb/t24/b1  ( .A(n559), .EN(n269), .Y(b[24]) );
  TBUFX2 \myram/m7/tb/t23/b1  ( .A(n558), .EN(n269), .Y(b[23]) );
  TBUFX2 \myram/m7/tb/t22/b1  ( .A(n557), .EN(n269), .Y(b[22]) );
  TBUFX2 \myram/m7/tb/t21/b1  ( .A(n556), .EN(n269), .Y(b[21]) );
  TBUFX2 \myram/m7/tb/t20/b1  ( .A(n555), .EN(n269), .Y(b[20]) );
  TBUFX2 \myram/m7/tb/t19/b1  ( .A(n554), .EN(n269), .Y(b[19]) );
  TBUFX2 \myram/m7/tb/t18/b1  ( .A(n553), .EN(n269), .Y(b[18]) );
  TBUFX2 \myram/m7/tb/t17/b1  ( .A(n552), .EN(n269), .Y(b[17]) );
  TBUFX2 \myram/m7/tb/t16/b1  ( .A(n551), .EN(n269), .Y(b[16]) );
  TBUFX2 \myram/m7/tb/t15/b1  ( .A(n550), .EN(n269), .Y(b[15]) );
  TBUFX2 \myram/m7/tb/t14/b1  ( .A(n549), .EN(n269), .Y(b[14]) );
  TBUFX2 \myram/m7/tb/t13/b1  ( .A(n548), .EN(n269), .Y(b[13]) );
  TBUFX2 \myram/m7/tb/t12/b1  ( .A(n547), .EN(n268), .Y(b[12]) );
  TBUFX2 \myram/m7/tb/t11/b1  ( .A(n546), .EN(n268), .Y(b[11]) );
  TBUFX2 \myram/m7/tb/t10/b1  ( .A(n545), .EN(n268), .Y(b[10]) );
  TBUFX2 \myram/m7/tb/t9/b1  ( .A(n544), .EN(n268), .Y(b[9]) );
  TBUFX2 \myram/m7/tb/t8/b1  ( .A(n543), .EN(n268), .Y(b[8]) );
  TBUFX2 \myram/m7/tb/t7/b1  ( .A(n542), .EN(n268), .Y(b[7]) );
  TBUFX2 \myram/m7/tb/t6/b1  ( .A(n541), .EN(n268), .Y(b[6]) );
  TBUFX2 \myram/m7/tb/t5/b1  ( .A(n540), .EN(n268), .Y(b[5]) );
  INVX1 \myram/m7/tb/t4/U1  ( .A(\myram/m7/dout[4] ), .Y(n571) );
  TBUFX2 \myram/m7/tb/t4/b1  ( .A(n571), .EN(n268), .Y(b[4]) );
  INVX1 \myram/m7/tb/t3/U1  ( .A(\myram/m7/dout[3] ), .Y(n570) );
  TBUFX2 \myram/m7/tb/t3/b1  ( .A(n570), .EN(n268), .Y(b[3]) );
  INVX1 \myram/m7/tb/t2/U1  ( .A(\myram/m7/dout[2] ), .Y(n569) );
  TBUFX2 \myram/m7/tb/t2/b1  ( .A(n569), .EN(n268), .Y(b[2]) );
  INVX1 \myram/m7/tb/t1/U1  ( .A(\myram/m7/dout[1] ), .Y(n568) );
  TBUFX2 \myram/m7/tb/t1/b1  ( .A(n568), .EN(n268), .Y(b[1]) );
  INVX1 \myram/m7/tb/t0/U1  ( .A(\myram/m7/dout[0] ), .Y(n567) );
  TBUFX2 \myram/m7/tb/t0/b1  ( .A(n567), .EN(n268), .Y(b[0]) );
  INVX1 \myram/m7/ta/t31/U1  ( .A(\myram/m7/dout[31] ), .Y(n566) );
  TBUFX2 \myram/m7/ta/t31/b1  ( .A(n566), .EN(\myram/sel_a[7] ), .Y(a[31]) );
  INVX1 \myram/m7/ta/t30/U1  ( .A(\myram/m7/dout[30] ), .Y(n565) );
  TBUFX2 \myram/m7/ta/t30/b1  ( .A(n565), .EN(\myram/sel_a[7] ), .Y(a[30]) );
  INVX1 \myram/m7/ta/t29/U1  ( .A(\myram/m7/dout[29] ), .Y(n564) );
  TBUFX2 \myram/m7/ta/t29/b1  ( .A(n564), .EN(\myram/sel_a[7] ), .Y(a[29]) );
  INVX1 \myram/m7/ta/t28/U1  ( .A(\myram/m7/dout[28] ), .Y(n563) );
  TBUFX2 \myram/m7/ta/t28/b1  ( .A(n563), .EN(\myram/sel_a[7] ), .Y(a[28]) );
  INVX1 \myram/m7/ta/t27/U1  ( .A(\myram/m7/dout[27] ), .Y(n562) );
  TBUFX2 \myram/m7/ta/t27/b1  ( .A(n562), .EN(\myram/sel_a[7] ), .Y(a[27]) );
  INVX1 \myram/m7/ta/t26/U1  ( .A(\myram/m7/dout[26] ), .Y(n561) );
  TBUFX2 \myram/m7/ta/t26/b1  ( .A(n561), .EN(\myram/sel_a[7] ), .Y(a[26]) );
  INVX1 \myram/m7/ta/t25/U1  ( .A(\myram/m7/dout[25] ), .Y(n560) );
  TBUFX2 \myram/m7/ta/t25/b1  ( .A(n560), .EN(\myram/sel_a[7] ), .Y(a[25]) );
  INVX1 \myram/m7/ta/t24/U1  ( .A(\myram/m7/dout[24] ), .Y(n559) );
  TBUFX2 \myram/m7/ta/t24/b1  ( .A(n559), .EN(\myram/sel_a[7] ), .Y(a[24]) );
  INVX1 \myram/m7/ta/t23/U1  ( .A(\myram/m7/dout[23] ), .Y(n558) );
  TBUFX2 \myram/m7/ta/t23/b1  ( .A(n558), .EN(\myram/sel_a[7] ), .Y(a[23]) );
  INVX1 \myram/m7/ta/t22/U1  ( .A(\myram/m7/dout[22] ), .Y(n557) );
  TBUFX2 \myram/m7/ta/t22/b1  ( .A(n557), .EN(\myram/sel_a[7] ), .Y(a[22]) );
  INVX1 \myram/m7/ta/t21/U1  ( .A(\myram/m7/dout[21] ), .Y(n556) );
  TBUFX2 \myram/m7/ta/t21/b1  ( .A(n556), .EN(\myram/sel_a[7] ), .Y(a[21]) );
  INVX1 \myram/m7/ta/t20/U1  ( .A(\myram/m7/dout[20] ), .Y(n555) );
  TBUFX2 \myram/m7/ta/t20/b1  ( .A(n555), .EN(\myram/sel_a[7] ), .Y(a[20]) );
  INVX1 \myram/m7/ta/t19/U1  ( .A(\myram/m7/dout[19] ), .Y(n554) );
  TBUFX2 \myram/m7/ta/t19/b1  ( .A(n554), .EN(\myram/sel_a[7] ), .Y(a[19]) );
  INVX1 \myram/m7/ta/t18/U1  ( .A(\myram/m7/dout[18] ), .Y(n553) );
  TBUFX2 \myram/m7/ta/t18/b1  ( .A(n553), .EN(\myram/sel_a[7] ), .Y(a[18]) );
  INVX1 \myram/m7/ta/t17/U1  ( .A(\myram/m7/dout[17] ), .Y(n552) );
  TBUFX2 \myram/m7/ta/t17/b1  ( .A(n552), .EN(\myram/sel_a[7] ), .Y(a[17]) );
  INVX1 \myram/m7/ta/t16/U1  ( .A(\myram/m7/dout[16] ), .Y(n551) );
  TBUFX2 \myram/m7/ta/t16/b1  ( .A(n551), .EN(\myram/sel_a[7] ), .Y(a[16]) );
  INVX1 \myram/m7/ta/t15/U1  ( .A(\myram/m7/dout[15] ), .Y(n550) );
  TBUFX2 \myram/m7/ta/t15/b1  ( .A(n550), .EN(\myram/sel_a[7] ), .Y(a[15]) );
  INVX1 \myram/m7/ta/t14/U1  ( .A(\myram/m7/dout[14] ), .Y(n549) );
  TBUFX2 \myram/m7/ta/t14/b1  ( .A(n549), .EN(\myram/sel_a[7] ), .Y(a[14]) );
  INVX1 \myram/m7/ta/t13/U1  ( .A(\myram/m7/dout[13] ), .Y(n548) );
  TBUFX2 \myram/m7/ta/t13/b1  ( .A(n548), .EN(n228), .Y(a[13]) );
  INVX1 \myram/m7/ta/t12/U1  ( .A(\myram/m7/dout[12] ), .Y(n547) );
  TBUFX2 \myram/m7/ta/t12/b1  ( .A(n547), .EN(n228), .Y(a[12]) );
  INVX1 \myram/m7/ta/t11/U1  ( .A(\myram/m7/dout[11] ), .Y(n546) );
  TBUFX2 \myram/m7/ta/t11/b1  ( .A(n546), .EN(n228), .Y(a[11]) );
  INVX1 \myram/m7/ta/t10/U1  ( .A(\myram/m7/dout[10] ), .Y(n545) );
  TBUFX2 \myram/m7/ta/t10/b1  ( .A(n545), .EN(n228), .Y(a[10]) );
  INVX1 \myram/m7/ta/t9/U1  ( .A(\myram/m7/dout[9] ), .Y(n544) );
  TBUFX2 \myram/m7/ta/t9/b1  ( .A(n544), .EN(n228), .Y(a[9]) );
  INVX1 \myram/m7/ta/t8/U1  ( .A(\myram/m7/dout[8] ), .Y(n543) );
  TBUFX2 \myram/m7/ta/t8/b1  ( .A(n543), .EN(n228), .Y(a[8]) );
  INVX1 \myram/m7/ta/t7/U1  ( .A(\myram/m7/dout[7] ), .Y(n542) );
  TBUFX2 \myram/m7/ta/t7/b1  ( .A(n542), .EN(n228), .Y(a[7]) );
  INVX1 \myram/m7/ta/t6/U1  ( .A(\myram/m7/dout[6] ), .Y(n541) );
  TBUFX2 \myram/m7/ta/t6/b1  ( .A(n541), .EN(n228), .Y(a[6]) );
  INVX1 \myram/m7/ta/t5/U1  ( .A(\myram/m7/dout[5] ), .Y(n540) );
  TBUFX2 \myram/m7/ta/t5/b1  ( .A(n540), .EN(n228), .Y(a[5]) );
  TBUFX2 \myram/m7/ta/t4/b1  ( .A(n571), .EN(n228), .Y(a[4]) );
  TBUFX2 \myram/m7/ta/t3/b1  ( .A(n570), .EN(n228), .Y(a[3]) );
  TBUFX2 \myram/m7/ta/t2/b1  ( .A(n569), .EN(n228), .Y(a[2]) );
  TBUFX2 \myram/m7/ta/t1/b1  ( .A(n568), .EN(n228), .Y(a[1]) );
  TBUFX2 \myram/m7/ta/t0/b1  ( .A(n567), .EN(n228), .Y(a[0]) );
  TBUFX2 \myram/m6/tb/t31/b1  ( .A(n534), .EN(n272), .Y(b[31]) );
  TBUFX2 \myram/m6/tb/t30/b1  ( .A(n533), .EN(n272), .Y(b[30]) );
  TBUFX2 \myram/m6/tb/t29/b1  ( .A(n532), .EN(n272), .Y(b[29]) );
  TBUFX2 \myram/m6/tb/t28/b1  ( .A(n531), .EN(n272), .Y(b[28]) );
  TBUFX2 \myram/m6/tb/t27/b1  ( .A(n530), .EN(n272), .Y(b[27]) );
  TBUFX2 \myram/m6/tb/t26/b1  ( .A(n529), .EN(n272), .Y(b[26]) );
  TBUFX2 \myram/m6/tb/t25/b1  ( .A(n528), .EN(n272), .Y(b[25]) );
  TBUFX2 \myram/m6/tb/t24/b1  ( .A(n527), .EN(n272), .Y(b[24]) );
  TBUFX2 \myram/m6/tb/t23/b1  ( .A(n526), .EN(n272), .Y(b[23]) );
  TBUFX2 \myram/m6/tb/t22/b1  ( .A(n525), .EN(n272), .Y(b[22]) );
  TBUFX2 \myram/m6/tb/t21/b1  ( .A(n524), .EN(n272), .Y(b[21]) );
  TBUFX2 \myram/m6/tb/t20/b1  ( .A(n523), .EN(n272), .Y(b[20]) );
  TBUFX2 \myram/m6/tb/t19/b1  ( .A(n522), .EN(n272), .Y(b[19]) );
  TBUFX2 \myram/m6/tb/t18/b1  ( .A(n521), .EN(n272), .Y(b[18]) );
  TBUFX2 \myram/m6/tb/t17/b1  ( .A(n520), .EN(n272), .Y(b[17]) );
  TBUFX2 \myram/m6/tb/t16/b1  ( .A(n519), .EN(n272), .Y(b[16]) );
  TBUFX2 \myram/m6/tb/t15/b1  ( .A(n518), .EN(n272), .Y(b[15]) );
  TBUFX2 \myram/m6/tb/t14/b1  ( .A(n517), .EN(n272), .Y(b[14]) );
  TBUFX2 \myram/m6/tb/t13/b1  ( .A(n516), .EN(n272), .Y(b[13]) );
  TBUFX2 \myram/m6/tb/t12/b1  ( .A(n515), .EN(n271), .Y(b[12]) );
  TBUFX2 \myram/m6/tb/t11/b1  ( .A(n514), .EN(n271), .Y(b[11]) );
  TBUFX2 \myram/m6/tb/t10/b1  ( .A(n513), .EN(n271), .Y(b[10]) );
  TBUFX2 \myram/m6/tb/t9/b1  ( .A(n512), .EN(n271), .Y(b[9]) );
  TBUFX2 \myram/m6/tb/t8/b1  ( .A(n511), .EN(n271), .Y(b[8]) );
  TBUFX2 \myram/m6/tb/t7/b1  ( .A(n510), .EN(n271), .Y(b[7]) );
  TBUFX2 \myram/m6/tb/t6/b1  ( .A(n509), .EN(n271), .Y(b[6]) );
  TBUFX2 \myram/m6/tb/t5/b1  ( .A(n508), .EN(n271), .Y(b[5]) );
  INVX1 \myram/m6/tb/t4/U1  ( .A(\myram/m6/dout[4] ), .Y(n539) );
  TBUFX2 \myram/m6/tb/t4/b1  ( .A(n539), .EN(n271), .Y(b[4]) );
  INVX1 \myram/m6/tb/t3/U1  ( .A(\myram/m6/dout[3] ), .Y(n538) );
  TBUFX2 \myram/m6/tb/t3/b1  ( .A(n538), .EN(n271), .Y(b[3]) );
  INVX1 \myram/m6/tb/t2/U1  ( .A(\myram/m6/dout[2] ), .Y(n537) );
  TBUFX2 \myram/m6/tb/t2/b1  ( .A(n537), .EN(n271), .Y(b[2]) );
  INVX1 \myram/m6/tb/t1/U1  ( .A(\myram/m6/dout[1] ), .Y(n536) );
  TBUFX2 \myram/m6/tb/t1/b1  ( .A(n536), .EN(n271), .Y(b[1]) );
  INVX1 \myram/m6/tb/t0/U1  ( .A(\myram/m6/dout[0] ), .Y(n535) );
  TBUFX2 \myram/m6/tb/t0/b1  ( .A(n535), .EN(n271), .Y(b[0]) );
  INVX1 \myram/m6/ta/t31/U1  ( .A(\myram/m6/dout[31] ), .Y(n534) );
  TBUFX2 \myram/m6/ta/t31/b1  ( .A(n534), .EN(\myram/sel_a[6] ), .Y(a[31]) );
  INVX1 \myram/m6/ta/t30/U1  ( .A(\myram/m6/dout[30] ), .Y(n533) );
  TBUFX2 \myram/m6/ta/t30/b1  ( .A(n533), .EN(\myram/sel_a[6] ), .Y(a[30]) );
  INVX1 \myram/m6/ta/t29/U1  ( .A(\myram/m6/dout[29] ), .Y(n532) );
  TBUFX2 \myram/m6/ta/t29/b1  ( .A(n532), .EN(\myram/sel_a[6] ), .Y(a[29]) );
  INVX1 \myram/m6/ta/t28/U1  ( .A(\myram/m6/dout[28] ), .Y(n531) );
  TBUFX2 \myram/m6/ta/t28/b1  ( .A(n531), .EN(\myram/sel_a[6] ), .Y(a[28]) );
  INVX1 \myram/m6/ta/t27/U1  ( .A(\myram/m6/dout[27] ), .Y(n530) );
  TBUFX2 \myram/m6/ta/t27/b1  ( .A(n530), .EN(\myram/sel_a[6] ), .Y(a[27]) );
  INVX1 \myram/m6/ta/t26/U1  ( .A(\myram/m6/dout[26] ), .Y(n529) );
  TBUFX2 \myram/m6/ta/t26/b1  ( .A(n529), .EN(\myram/sel_a[6] ), .Y(a[26]) );
  INVX1 \myram/m6/ta/t25/U1  ( .A(\myram/m6/dout[25] ), .Y(n528) );
  TBUFX2 \myram/m6/ta/t25/b1  ( .A(n528), .EN(\myram/sel_a[6] ), .Y(a[25]) );
  INVX1 \myram/m6/ta/t24/U1  ( .A(\myram/m6/dout[24] ), .Y(n527) );
  TBUFX2 \myram/m6/ta/t24/b1  ( .A(n527), .EN(\myram/sel_a[6] ), .Y(a[24]) );
  INVX1 \myram/m6/ta/t23/U1  ( .A(\myram/m6/dout[23] ), .Y(n526) );
  TBUFX2 \myram/m6/ta/t23/b1  ( .A(n526), .EN(\myram/sel_a[6] ), .Y(a[23]) );
  INVX1 \myram/m6/ta/t22/U1  ( .A(\myram/m6/dout[22] ), .Y(n525) );
  TBUFX2 \myram/m6/ta/t22/b1  ( .A(n525), .EN(\myram/sel_a[6] ), .Y(a[22]) );
  INVX1 \myram/m6/ta/t21/U1  ( .A(\myram/m6/dout[21] ), .Y(n524) );
  TBUFX2 \myram/m6/ta/t21/b1  ( .A(n524), .EN(\myram/sel_a[6] ), .Y(a[21]) );
  INVX1 \myram/m6/ta/t20/U1  ( .A(\myram/m6/dout[20] ), .Y(n523) );
  TBUFX2 \myram/m6/ta/t20/b1  ( .A(n523), .EN(\myram/sel_a[6] ), .Y(a[20]) );
  INVX1 \myram/m6/ta/t19/U1  ( .A(\myram/m6/dout[19] ), .Y(n522) );
  TBUFX2 \myram/m6/ta/t19/b1  ( .A(n522), .EN(\myram/sel_a[6] ), .Y(a[19]) );
  INVX1 \myram/m6/ta/t18/U1  ( .A(\myram/m6/dout[18] ), .Y(n521) );
  TBUFX2 \myram/m6/ta/t18/b1  ( .A(n521), .EN(\myram/sel_a[6] ), .Y(a[18]) );
  INVX1 \myram/m6/ta/t17/U1  ( .A(\myram/m6/dout[17] ), .Y(n520) );
  TBUFX2 \myram/m6/ta/t17/b1  ( .A(n520), .EN(\myram/sel_a[6] ), .Y(a[17]) );
  INVX1 \myram/m6/ta/t16/U1  ( .A(\myram/m6/dout[16] ), .Y(n519) );
  TBUFX2 \myram/m6/ta/t16/b1  ( .A(n519), .EN(\myram/sel_a[6] ), .Y(a[16]) );
  INVX1 \myram/m6/ta/t15/U1  ( .A(\myram/m6/dout[15] ), .Y(n518) );
  TBUFX2 \myram/m6/ta/t15/b1  ( .A(n518), .EN(\myram/sel_a[6] ), .Y(a[15]) );
  INVX1 \myram/m6/ta/t14/U1  ( .A(\myram/m6/dout[14] ), .Y(n517) );
  TBUFX2 \myram/m6/ta/t14/b1  ( .A(n517), .EN(\myram/sel_a[6] ), .Y(a[14]) );
  INVX1 \myram/m6/ta/t13/U1  ( .A(\myram/m6/dout[13] ), .Y(n516) );
  TBUFX2 \myram/m6/ta/t13/b1  ( .A(n516), .EN(n230), .Y(a[13]) );
  INVX1 \myram/m6/ta/t12/U1  ( .A(\myram/m6/dout[12] ), .Y(n515) );
  TBUFX2 \myram/m6/ta/t12/b1  ( .A(n515), .EN(n230), .Y(a[12]) );
  INVX1 \myram/m6/ta/t11/U1  ( .A(\myram/m6/dout[11] ), .Y(n514) );
  TBUFX2 \myram/m6/ta/t11/b1  ( .A(n514), .EN(n230), .Y(a[11]) );
  INVX1 \myram/m6/ta/t10/U1  ( .A(\myram/m6/dout[10] ), .Y(n513) );
  TBUFX2 \myram/m6/ta/t10/b1  ( .A(n513), .EN(n230), .Y(a[10]) );
  INVX1 \myram/m6/ta/t9/U1  ( .A(\myram/m6/dout[9] ), .Y(n512) );
  TBUFX2 \myram/m6/ta/t9/b1  ( .A(n512), .EN(n230), .Y(a[9]) );
  INVX1 \myram/m6/ta/t8/U1  ( .A(\myram/m6/dout[8] ), .Y(n511) );
  TBUFX2 \myram/m6/ta/t8/b1  ( .A(n511), .EN(n230), .Y(a[8]) );
  INVX1 \myram/m6/ta/t7/U1  ( .A(\myram/m6/dout[7] ), .Y(n510) );
  TBUFX2 \myram/m6/ta/t7/b1  ( .A(n510), .EN(n230), .Y(a[7]) );
  INVX1 \myram/m6/ta/t6/U1  ( .A(\myram/m6/dout[6] ), .Y(n509) );
  TBUFX2 \myram/m6/ta/t6/b1  ( .A(n509), .EN(n230), .Y(a[6]) );
  INVX1 \myram/m6/ta/t5/U1  ( .A(\myram/m6/dout[5] ), .Y(n508) );
  TBUFX2 \myram/m6/ta/t5/b1  ( .A(n508), .EN(n230), .Y(a[5]) );
  TBUFX2 \myram/m6/ta/t4/b1  ( .A(n539), .EN(n230), .Y(a[4]) );
  TBUFX2 \myram/m6/ta/t3/b1  ( .A(n538), .EN(n230), .Y(a[3]) );
  TBUFX2 \myram/m6/ta/t2/b1  ( .A(n537), .EN(n230), .Y(a[2]) );
  TBUFX2 \myram/m6/ta/t1/b1  ( .A(n536), .EN(n230), .Y(a[1]) );
  TBUFX2 \myram/m6/ta/t0/b1  ( .A(n535), .EN(n230), .Y(a[0]) );
  TBUFX2 \myram/m5/tb/t31/b1  ( .A(n502), .EN(n275), .Y(b[31]) );
  TBUFX2 \myram/m5/tb/t30/b1  ( .A(n501), .EN(n275), .Y(b[30]) );
  TBUFX2 \myram/m5/tb/t29/b1  ( .A(n500), .EN(n275), .Y(b[29]) );
  TBUFX2 \myram/m5/tb/t28/b1  ( .A(n499), .EN(n275), .Y(b[28]) );
  TBUFX2 \myram/m5/tb/t27/b1  ( .A(n498), .EN(n275), .Y(b[27]) );
  TBUFX2 \myram/m5/tb/t26/b1  ( .A(n497), .EN(n275), .Y(b[26]) );
  TBUFX2 \myram/m5/tb/t25/b1  ( .A(n496), .EN(n275), .Y(b[25]) );
  TBUFX2 \myram/m5/tb/t24/b1  ( .A(n495), .EN(n275), .Y(b[24]) );
  TBUFX2 \myram/m5/tb/t23/b1  ( .A(n494), .EN(n275), .Y(b[23]) );
  TBUFX2 \myram/m5/tb/t22/b1  ( .A(n493), .EN(n275), .Y(b[22]) );
  TBUFX2 \myram/m5/tb/t21/b1  ( .A(n492), .EN(n275), .Y(b[21]) );
  TBUFX2 \myram/m5/tb/t20/b1  ( .A(n491), .EN(n275), .Y(b[20]) );
  TBUFX2 \myram/m5/tb/t19/b1  ( .A(n490), .EN(n275), .Y(b[19]) );
  TBUFX2 \myram/m5/tb/t18/b1  ( .A(n489), .EN(n275), .Y(b[18]) );
  TBUFX2 \myram/m5/tb/t17/b1  ( .A(n488), .EN(n275), .Y(b[17]) );
  TBUFX2 \myram/m5/tb/t16/b1  ( .A(n487), .EN(n275), .Y(b[16]) );
  TBUFX2 \myram/m5/tb/t15/b1  ( .A(n486), .EN(n275), .Y(b[15]) );
  TBUFX2 \myram/m5/tb/t14/b1  ( .A(n485), .EN(n275), .Y(b[14]) );
  TBUFX2 \myram/m5/tb/t13/b1  ( .A(n484), .EN(n275), .Y(b[13]) );
  TBUFX2 \myram/m5/tb/t12/b1  ( .A(n483), .EN(n274), .Y(b[12]) );
  TBUFX2 \myram/m5/tb/t11/b1  ( .A(n482), .EN(n274), .Y(b[11]) );
  TBUFX2 \myram/m5/tb/t10/b1  ( .A(n481), .EN(n274), .Y(b[10]) );
  TBUFX2 \myram/m5/tb/t9/b1  ( .A(n480), .EN(n274), .Y(b[9]) );
  TBUFX2 \myram/m5/tb/t8/b1  ( .A(n479), .EN(n274), .Y(b[8]) );
  TBUFX2 \myram/m5/tb/t7/b1  ( .A(n478), .EN(n274), .Y(b[7]) );
  TBUFX2 \myram/m5/tb/t6/b1  ( .A(n477), .EN(n274), .Y(b[6]) );
  TBUFX2 \myram/m5/tb/t5/b1  ( .A(n476), .EN(n274), .Y(b[5]) );
  INVX1 \myram/m5/tb/t4/U1  ( .A(\myram/m5/dout[4] ), .Y(n507) );
  TBUFX2 \myram/m5/tb/t4/b1  ( .A(n507), .EN(n274), .Y(b[4]) );
  INVX1 \myram/m5/tb/t3/U1  ( .A(\myram/m5/dout[3] ), .Y(n506) );
  TBUFX2 \myram/m5/tb/t3/b1  ( .A(n506), .EN(n274), .Y(b[3]) );
  INVX1 \myram/m5/tb/t2/U1  ( .A(\myram/m5/dout[2] ), .Y(n505) );
  TBUFX2 \myram/m5/tb/t2/b1  ( .A(n505), .EN(n274), .Y(b[2]) );
  INVX1 \myram/m5/tb/t1/U1  ( .A(\myram/m5/dout[1] ), .Y(n504) );
  TBUFX2 \myram/m5/tb/t1/b1  ( .A(n504), .EN(n274), .Y(b[1]) );
  INVX1 \myram/m5/tb/t0/U1  ( .A(\myram/m5/dout[0] ), .Y(n503) );
  TBUFX2 \myram/m5/tb/t0/b1  ( .A(n503), .EN(n274), .Y(b[0]) );
  INVX1 \myram/m5/ta/t31/U1  ( .A(\myram/m5/dout[31] ), .Y(n502) );
  TBUFX2 \myram/m5/ta/t31/b1  ( .A(n502), .EN(\myram/sel_a[5] ), .Y(a[31]) );
  INVX1 \myram/m5/ta/t30/U1  ( .A(\myram/m5/dout[30] ), .Y(n501) );
  TBUFX2 \myram/m5/ta/t30/b1  ( .A(n501), .EN(\myram/sel_a[5] ), .Y(a[30]) );
  INVX1 \myram/m5/ta/t29/U1  ( .A(\myram/m5/dout[29] ), .Y(n500) );
  TBUFX2 \myram/m5/ta/t29/b1  ( .A(n500), .EN(\myram/sel_a[5] ), .Y(a[29]) );
  INVX1 \myram/m5/ta/t28/U1  ( .A(\myram/m5/dout[28] ), .Y(n499) );
  TBUFX2 \myram/m5/ta/t28/b1  ( .A(n499), .EN(\myram/sel_a[5] ), .Y(a[28]) );
  INVX1 \myram/m5/ta/t27/U1  ( .A(\myram/m5/dout[27] ), .Y(n498) );
  TBUFX2 \myram/m5/ta/t27/b1  ( .A(n498), .EN(\myram/sel_a[5] ), .Y(a[27]) );
  INVX1 \myram/m5/ta/t26/U1  ( .A(\myram/m5/dout[26] ), .Y(n497) );
  TBUFX2 \myram/m5/ta/t26/b1  ( .A(n497), .EN(\myram/sel_a[5] ), .Y(a[26]) );
  INVX1 \myram/m5/ta/t25/U1  ( .A(\myram/m5/dout[25] ), .Y(n496) );
  TBUFX2 \myram/m5/ta/t25/b1  ( .A(n496), .EN(\myram/sel_a[5] ), .Y(a[25]) );
  INVX1 \myram/m5/ta/t24/U1  ( .A(\myram/m5/dout[24] ), .Y(n495) );
  TBUFX2 \myram/m5/ta/t24/b1  ( .A(n495), .EN(\myram/sel_a[5] ), .Y(a[24]) );
  INVX1 \myram/m5/ta/t23/U1  ( .A(\myram/m5/dout[23] ), .Y(n494) );
  TBUFX2 \myram/m5/ta/t23/b1  ( .A(n494), .EN(\myram/sel_a[5] ), .Y(a[23]) );
  INVX1 \myram/m5/ta/t22/U1  ( .A(\myram/m5/dout[22] ), .Y(n493) );
  TBUFX2 \myram/m5/ta/t22/b1  ( .A(n493), .EN(\myram/sel_a[5] ), .Y(a[22]) );
  INVX1 \myram/m5/ta/t21/U1  ( .A(\myram/m5/dout[21] ), .Y(n492) );
  TBUFX2 \myram/m5/ta/t21/b1  ( .A(n492), .EN(\myram/sel_a[5] ), .Y(a[21]) );
  INVX1 \myram/m5/ta/t20/U1  ( .A(\myram/m5/dout[20] ), .Y(n491) );
  TBUFX2 \myram/m5/ta/t20/b1  ( .A(n491), .EN(\myram/sel_a[5] ), .Y(a[20]) );
  INVX1 \myram/m5/ta/t19/U1  ( .A(\myram/m5/dout[19] ), .Y(n490) );
  TBUFX2 \myram/m5/ta/t19/b1  ( .A(n490), .EN(\myram/sel_a[5] ), .Y(a[19]) );
  INVX1 \myram/m5/ta/t18/U1  ( .A(\myram/m5/dout[18] ), .Y(n489) );
  TBUFX2 \myram/m5/ta/t18/b1  ( .A(n489), .EN(\myram/sel_a[5] ), .Y(a[18]) );
  INVX1 \myram/m5/ta/t17/U1  ( .A(\myram/m5/dout[17] ), .Y(n488) );
  TBUFX2 \myram/m5/ta/t17/b1  ( .A(n488), .EN(\myram/sel_a[5] ), .Y(a[17]) );
  INVX1 \myram/m5/ta/t16/U1  ( .A(\myram/m5/dout[16] ), .Y(n487) );
  TBUFX2 \myram/m5/ta/t16/b1  ( .A(n487), .EN(\myram/sel_a[5] ), .Y(a[16]) );
  INVX1 \myram/m5/ta/t15/U1  ( .A(\myram/m5/dout[15] ), .Y(n486) );
  TBUFX2 \myram/m5/ta/t15/b1  ( .A(n486), .EN(\myram/sel_a[5] ), .Y(a[15]) );
  INVX1 \myram/m5/ta/t14/U1  ( .A(\myram/m5/dout[14] ), .Y(n485) );
  TBUFX2 \myram/m5/ta/t14/b1  ( .A(n485), .EN(\myram/sel_a[5] ), .Y(a[14]) );
  INVX1 \myram/m5/ta/t13/U1  ( .A(\myram/m5/dout[13] ), .Y(n484) );
  TBUFX2 \myram/m5/ta/t13/b1  ( .A(n484), .EN(n232), .Y(a[13]) );
  INVX1 \myram/m5/ta/t12/U1  ( .A(\myram/m5/dout[12] ), .Y(n483) );
  TBUFX2 \myram/m5/ta/t12/b1  ( .A(n483), .EN(n232), .Y(a[12]) );
  INVX1 \myram/m5/ta/t11/U1  ( .A(\myram/m5/dout[11] ), .Y(n482) );
  TBUFX2 \myram/m5/ta/t11/b1  ( .A(n482), .EN(n232), .Y(a[11]) );
  INVX1 \myram/m5/ta/t10/U1  ( .A(\myram/m5/dout[10] ), .Y(n481) );
  TBUFX2 \myram/m5/ta/t10/b1  ( .A(n481), .EN(n232), .Y(a[10]) );
  INVX1 \myram/m5/ta/t9/U1  ( .A(\myram/m5/dout[9] ), .Y(n480) );
  TBUFX2 \myram/m5/ta/t9/b1  ( .A(n480), .EN(n232), .Y(a[9]) );
  INVX1 \myram/m5/ta/t8/U1  ( .A(\myram/m5/dout[8] ), .Y(n479) );
  TBUFX2 \myram/m5/ta/t8/b1  ( .A(n479), .EN(n232), .Y(a[8]) );
  INVX1 \myram/m5/ta/t7/U1  ( .A(\myram/m5/dout[7] ), .Y(n478) );
  TBUFX2 \myram/m5/ta/t7/b1  ( .A(n478), .EN(n232), .Y(a[7]) );
  INVX1 \myram/m5/ta/t6/U1  ( .A(\myram/m5/dout[6] ), .Y(n477) );
  TBUFX2 \myram/m5/ta/t6/b1  ( .A(n477), .EN(n232), .Y(a[6]) );
  INVX1 \myram/m5/ta/t5/U1  ( .A(\myram/m5/dout[5] ), .Y(n476) );
  TBUFX2 \myram/m5/ta/t5/b1  ( .A(n476), .EN(n232), .Y(a[5]) );
  TBUFX2 \myram/m5/ta/t4/b1  ( .A(n507), .EN(n232), .Y(a[4]) );
  TBUFX2 \myram/m5/ta/t3/b1  ( .A(n506), .EN(n232), .Y(a[3]) );
  TBUFX2 \myram/m5/ta/t2/b1  ( .A(n505), .EN(n232), .Y(a[2]) );
  TBUFX2 \myram/m5/ta/t1/b1  ( .A(n504), .EN(n232), .Y(a[1]) );
  TBUFX2 \myram/m5/ta/t0/b1  ( .A(n503), .EN(n232), .Y(a[0]) );
  TBUFX2 \myram/m4/tb/t31/b1  ( .A(n470), .EN(n278), .Y(b[31]) );
  TBUFX2 \myram/m4/tb/t30/b1  ( .A(n469), .EN(n278), .Y(b[30]) );
  TBUFX2 \myram/m4/tb/t29/b1  ( .A(n468), .EN(n278), .Y(b[29]) );
  TBUFX2 \myram/m4/tb/t28/b1  ( .A(n467), .EN(n278), .Y(b[28]) );
  TBUFX2 \myram/m4/tb/t27/b1  ( .A(n466), .EN(n278), .Y(b[27]) );
  TBUFX2 \myram/m4/tb/t26/b1  ( .A(n465), .EN(n278), .Y(b[26]) );
  TBUFX2 \myram/m4/tb/t25/b1  ( .A(n464), .EN(n278), .Y(b[25]) );
  TBUFX2 \myram/m4/tb/t24/b1  ( .A(n463), .EN(n278), .Y(b[24]) );
  TBUFX2 \myram/m4/tb/t23/b1  ( .A(n462), .EN(n278), .Y(b[23]) );
  TBUFX2 \myram/m4/tb/t22/b1  ( .A(n461), .EN(n278), .Y(b[22]) );
  TBUFX2 \myram/m4/tb/t21/b1  ( .A(n460), .EN(n278), .Y(b[21]) );
  TBUFX2 \myram/m4/tb/t20/b1  ( .A(n459), .EN(n278), .Y(b[20]) );
  TBUFX2 \myram/m4/tb/t19/b1  ( .A(n458), .EN(n278), .Y(b[19]) );
  TBUFX2 \myram/m4/tb/t18/b1  ( .A(n457), .EN(n278), .Y(b[18]) );
  TBUFX2 \myram/m4/tb/t17/b1  ( .A(n456), .EN(n278), .Y(b[17]) );
  TBUFX2 \myram/m4/tb/t16/b1  ( .A(n455), .EN(n278), .Y(b[16]) );
  TBUFX2 \myram/m4/tb/t15/b1  ( .A(n454), .EN(n278), .Y(b[15]) );
  TBUFX2 \myram/m4/tb/t14/b1  ( .A(n453), .EN(n278), .Y(b[14]) );
  TBUFX2 \myram/m4/tb/t13/b1  ( .A(n452), .EN(n278), .Y(b[13]) );
  TBUFX2 \myram/m4/tb/t12/b1  ( .A(n451), .EN(n277), .Y(b[12]) );
  TBUFX2 \myram/m4/tb/t11/b1  ( .A(n450), .EN(n277), .Y(b[11]) );
  TBUFX2 \myram/m4/tb/t10/b1  ( .A(n449), .EN(n277), .Y(b[10]) );
  TBUFX2 \myram/m4/tb/t9/b1  ( .A(n448), .EN(n277), .Y(b[9]) );
  TBUFX2 \myram/m4/tb/t8/b1  ( .A(n447), .EN(n277), .Y(b[8]) );
  TBUFX2 \myram/m4/tb/t7/b1  ( .A(n446), .EN(n277), .Y(b[7]) );
  TBUFX2 \myram/m4/tb/t6/b1  ( .A(n445), .EN(n277), .Y(b[6]) );
  TBUFX2 \myram/m4/tb/t5/b1  ( .A(n444), .EN(n277), .Y(b[5]) );
  INVX1 \myram/m4/tb/t4/U1  ( .A(\myram/m4/dout[4] ), .Y(n475) );
  TBUFX2 \myram/m4/tb/t4/b1  ( .A(n475), .EN(n277), .Y(b[4]) );
  INVX1 \myram/m4/tb/t3/U1  ( .A(\myram/m4/dout[3] ), .Y(n474) );
  TBUFX2 \myram/m4/tb/t3/b1  ( .A(n474), .EN(n277), .Y(b[3]) );
  INVX1 \myram/m4/tb/t2/U1  ( .A(\myram/m4/dout[2] ), .Y(n473) );
  TBUFX2 \myram/m4/tb/t2/b1  ( .A(n473), .EN(n277), .Y(b[2]) );
  INVX1 \myram/m4/tb/t1/U1  ( .A(\myram/m4/dout[1] ), .Y(n472) );
  TBUFX2 \myram/m4/tb/t1/b1  ( .A(n472), .EN(n277), .Y(b[1]) );
  INVX1 \myram/m4/tb/t0/U1  ( .A(\myram/m4/dout[0] ), .Y(n471) );
  TBUFX2 \myram/m4/tb/t0/b1  ( .A(n471), .EN(n277), .Y(b[0]) );
  INVX1 \myram/m4/ta/t31/U1  ( .A(\myram/m4/dout[31] ), .Y(n470) );
  TBUFX2 \myram/m4/ta/t31/b1  ( .A(n470), .EN(\myram/sel_a[4] ), .Y(a[31]) );
  INVX1 \myram/m4/ta/t30/U1  ( .A(\myram/m4/dout[30] ), .Y(n469) );
  TBUFX2 \myram/m4/ta/t30/b1  ( .A(n469), .EN(\myram/sel_a[4] ), .Y(a[30]) );
  INVX1 \myram/m4/ta/t29/U1  ( .A(\myram/m4/dout[29] ), .Y(n468) );
  TBUFX2 \myram/m4/ta/t29/b1  ( .A(n468), .EN(\myram/sel_a[4] ), .Y(a[29]) );
  INVX1 \myram/m4/ta/t28/U1  ( .A(\myram/m4/dout[28] ), .Y(n467) );
  TBUFX2 \myram/m4/ta/t28/b1  ( .A(n467), .EN(\myram/sel_a[4] ), .Y(a[28]) );
  INVX1 \myram/m4/ta/t27/U1  ( .A(\myram/m4/dout[27] ), .Y(n466) );
  TBUFX2 \myram/m4/ta/t27/b1  ( .A(n466), .EN(\myram/sel_a[4] ), .Y(a[27]) );
  INVX1 \myram/m4/ta/t26/U1  ( .A(\myram/m4/dout[26] ), .Y(n465) );
  TBUFX2 \myram/m4/ta/t26/b1  ( .A(n465), .EN(\myram/sel_a[4] ), .Y(a[26]) );
  INVX1 \myram/m4/ta/t25/U1  ( .A(\myram/m4/dout[25] ), .Y(n464) );
  TBUFX2 \myram/m4/ta/t25/b1  ( .A(n464), .EN(\myram/sel_a[4] ), .Y(a[25]) );
  INVX1 \myram/m4/ta/t24/U1  ( .A(\myram/m4/dout[24] ), .Y(n463) );
  TBUFX2 \myram/m4/ta/t24/b1  ( .A(n463), .EN(\myram/sel_a[4] ), .Y(a[24]) );
  INVX1 \myram/m4/ta/t23/U1  ( .A(\myram/m4/dout[23] ), .Y(n462) );
  TBUFX2 \myram/m4/ta/t23/b1  ( .A(n462), .EN(\myram/sel_a[4] ), .Y(a[23]) );
  INVX1 \myram/m4/ta/t22/U1  ( .A(\myram/m4/dout[22] ), .Y(n461) );
  TBUFX2 \myram/m4/ta/t22/b1  ( .A(n461), .EN(\myram/sel_a[4] ), .Y(a[22]) );
  INVX1 \myram/m4/ta/t21/U1  ( .A(\myram/m4/dout[21] ), .Y(n460) );
  TBUFX2 \myram/m4/ta/t21/b1  ( .A(n460), .EN(\myram/sel_a[4] ), .Y(a[21]) );
  INVX1 \myram/m4/ta/t20/U1  ( .A(\myram/m4/dout[20] ), .Y(n459) );
  TBUFX2 \myram/m4/ta/t20/b1  ( .A(n459), .EN(\myram/sel_a[4] ), .Y(a[20]) );
  INVX1 \myram/m4/ta/t19/U1  ( .A(\myram/m4/dout[19] ), .Y(n458) );
  TBUFX2 \myram/m4/ta/t19/b1  ( .A(n458), .EN(\myram/sel_a[4] ), .Y(a[19]) );
  INVX1 \myram/m4/ta/t18/U1  ( .A(\myram/m4/dout[18] ), .Y(n457) );
  TBUFX2 \myram/m4/ta/t18/b1  ( .A(n457), .EN(\myram/sel_a[4] ), .Y(a[18]) );
  INVX1 \myram/m4/ta/t17/U1  ( .A(\myram/m4/dout[17] ), .Y(n456) );
  TBUFX2 \myram/m4/ta/t17/b1  ( .A(n456), .EN(\myram/sel_a[4] ), .Y(a[17]) );
  INVX1 \myram/m4/ta/t16/U1  ( .A(\myram/m4/dout[16] ), .Y(n455) );
  TBUFX2 \myram/m4/ta/t16/b1  ( .A(n455), .EN(\myram/sel_a[4] ), .Y(a[16]) );
  INVX1 \myram/m4/ta/t15/U1  ( .A(\myram/m4/dout[15] ), .Y(n454) );
  TBUFX2 \myram/m4/ta/t15/b1  ( .A(n454), .EN(\myram/sel_a[4] ), .Y(a[15]) );
  INVX1 \myram/m4/ta/t14/U1  ( .A(\myram/m4/dout[14] ), .Y(n453) );
  TBUFX2 \myram/m4/ta/t14/b1  ( .A(n453), .EN(\myram/sel_a[4] ), .Y(a[14]) );
  INVX1 \myram/m4/ta/t13/U1  ( .A(\myram/m4/dout[13] ), .Y(n452) );
  TBUFX2 \myram/m4/ta/t13/b1  ( .A(n452), .EN(n234), .Y(a[13]) );
  INVX1 \myram/m4/ta/t12/U1  ( .A(\myram/m4/dout[12] ), .Y(n451) );
  TBUFX2 \myram/m4/ta/t12/b1  ( .A(n451), .EN(n234), .Y(a[12]) );
  INVX1 \myram/m4/ta/t11/U1  ( .A(\myram/m4/dout[11] ), .Y(n450) );
  TBUFX2 \myram/m4/ta/t11/b1  ( .A(n450), .EN(n234), .Y(a[11]) );
  INVX1 \myram/m4/ta/t10/U1  ( .A(\myram/m4/dout[10] ), .Y(n449) );
  TBUFX2 \myram/m4/ta/t10/b1  ( .A(n449), .EN(n234), .Y(a[10]) );
  INVX1 \myram/m4/ta/t9/U1  ( .A(\myram/m4/dout[9] ), .Y(n448) );
  TBUFX2 \myram/m4/ta/t9/b1  ( .A(n448), .EN(n234), .Y(a[9]) );
  INVX1 \myram/m4/ta/t8/U1  ( .A(\myram/m4/dout[8] ), .Y(n447) );
  TBUFX2 \myram/m4/ta/t8/b1  ( .A(n447), .EN(n234), .Y(a[8]) );
  INVX1 \myram/m4/ta/t7/U1  ( .A(\myram/m4/dout[7] ), .Y(n446) );
  TBUFX2 \myram/m4/ta/t7/b1  ( .A(n446), .EN(n234), .Y(a[7]) );
  INVX1 \myram/m4/ta/t6/U1  ( .A(\myram/m4/dout[6] ), .Y(n445) );
  TBUFX2 \myram/m4/ta/t6/b1  ( .A(n445), .EN(n234), .Y(a[6]) );
  INVX1 \myram/m4/ta/t5/U1  ( .A(\myram/m4/dout[5] ), .Y(n444) );
  TBUFX2 \myram/m4/ta/t5/b1  ( .A(n444), .EN(n234), .Y(a[5]) );
  TBUFX2 \myram/m4/ta/t4/b1  ( .A(n475), .EN(n234), .Y(a[4]) );
  TBUFX2 \myram/m4/ta/t3/b1  ( .A(n474), .EN(n234), .Y(a[3]) );
  TBUFX2 \myram/m4/ta/t2/b1  ( .A(n473), .EN(n234), .Y(a[2]) );
  TBUFX2 \myram/m4/ta/t1/b1  ( .A(n472), .EN(n234), .Y(a[1]) );
  TBUFX2 \myram/m4/ta/t0/b1  ( .A(n471), .EN(n234), .Y(a[0]) );
  TBUFX2 \myram/m3/tb/t31/b1  ( .A(n438), .EN(n281), .Y(b[31]) );
  TBUFX2 \myram/m3/tb/t30/b1  ( .A(n437), .EN(n281), .Y(b[30]) );
  TBUFX2 \myram/m3/tb/t29/b1  ( .A(n436), .EN(n281), .Y(b[29]) );
  TBUFX2 \myram/m3/tb/t28/b1  ( .A(n435), .EN(n281), .Y(b[28]) );
  TBUFX2 \myram/m3/tb/t27/b1  ( .A(n434), .EN(n281), .Y(b[27]) );
  TBUFX2 \myram/m3/tb/t26/b1  ( .A(n433), .EN(n281), .Y(b[26]) );
  TBUFX2 \myram/m3/tb/t25/b1  ( .A(n432), .EN(n281), .Y(b[25]) );
  TBUFX2 \myram/m3/tb/t24/b1  ( .A(n431), .EN(n281), .Y(b[24]) );
  TBUFX2 \myram/m3/tb/t23/b1  ( .A(n430), .EN(n281), .Y(b[23]) );
  TBUFX2 \myram/m3/tb/t22/b1  ( .A(n429), .EN(n281), .Y(b[22]) );
  TBUFX2 \myram/m3/tb/t21/b1  ( .A(n428), .EN(n281), .Y(b[21]) );
  TBUFX2 \myram/m3/tb/t20/b1  ( .A(n427), .EN(n281), .Y(b[20]) );
  TBUFX2 \myram/m3/tb/t19/b1  ( .A(n426), .EN(n281), .Y(b[19]) );
  TBUFX2 \myram/m3/tb/t18/b1  ( .A(n425), .EN(n281), .Y(b[18]) );
  TBUFX2 \myram/m3/tb/t17/b1  ( .A(n424), .EN(n281), .Y(b[17]) );
  TBUFX2 \myram/m3/tb/t16/b1  ( .A(n423), .EN(n281), .Y(b[16]) );
  TBUFX2 \myram/m3/tb/t15/b1  ( .A(n422), .EN(n281), .Y(b[15]) );
  TBUFX2 \myram/m3/tb/t14/b1  ( .A(n421), .EN(n281), .Y(b[14]) );
  TBUFX2 \myram/m3/tb/t13/b1  ( .A(n420), .EN(n281), .Y(b[13]) );
  TBUFX2 \myram/m3/tb/t12/b1  ( .A(n419), .EN(n280), .Y(b[12]) );
  TBUFX2 \myram/m3/tb/t11/b1  ( .A(n418), .EN(n280), .Y(b[11]) );
  TBUFX2 \myram/m3/tb/t10/b1  ( .A(n417), .EN(n280), .Y(b[10]) );
  TBUFX2 \myram/m3/tb/t9/b1  ( .A(n416), .EN(n280), .Y(b[9]) );
  TBUFX2 \myram/m3/tb/t8/b1  ( .A(n415), .EN(n280), .Y(b[8]) );
  TBUFX2 \myram/m3/tb/t7/b1  ( .A(n414), .EN(n280), .Y(b[7]) );
  TBUFX2 \myram/m3/tb/t6/b1  ( .A(n413), .EN(n280), .Y(b[6]) );
  TBUFX2 \myram/m3/tb/t5/b1  ( .A(n412), .EN(n280), .Y(b[5]) );
  INVX1 \myram/m3/tb/t4/U1  ( .A(\myram/m3/dout[4] ), .Y(n443) );
  TBUFX2 \myram/m3/tb/t4/b1  ( .A(n443), .EN(n280), .Y(b[4]) );
  INVX1 \myram/m3/tb/t3/U1  ( .A(\myram/m3/dout[3] ), .Y(n442) );
  TBUFX2 \myram/m3/tb/t3/b1  ( .A(n442), .EN(n280), .Y(b[3]) );
  INVX1 \myram/m3/tb/t2/U1  ( .A(\myram/m3/dout[2] ), .Y(n441) );
  TBUFX2 \myram/m3/tb/t2/b1  ( .A(n441), .EN(n280), .Y(b[2]) );
  INVX1 \myram/m3/tb/t1/U1  ( .A(\myram/m3/dout[1] ), .Y(n440) );
  TBUFX2 \myram/m3/tb/t1/b1  ( .A(n440), .EN(n280), .Y(b[1]) );
  INVX1 \myram/m3/tb/t0/U1  ( .A(\myram/m3/dout[0] ), .Y(n439) );
  TBUFX2 \myram/m3/tb/t0/b1  ( .A(n439), .EN(n280), .Y(b[0]) );
  INVX1 \myram/m3/ta/t31/U1  ( .A(\myram/m3/dout[31] ), .Y(n438) );
  TBUFX2 \myram/m3/ta/t31/b1  ( .A(n438), .EN(\myram/sel_a[3] ), .Y(a[31]) );
  INVX1 \myram/m3/ta/t30/U1  ( .A(\myram/m3/dout[30] ), .Y(n437) );
  TBUFX2 \myram/m3/ta/t30/b1  ( .A(n437), .EN(\myram/sel_a[3] ), .Y(a[30]) );
  INVX1 \myram/m3/ta/t29/U1  ( .A(\myram/m3/dout[29] ), .Y(n436) );
  TBUFX2 \myram/m3/ta/t29/b1  ( .A(n436), .EN(\myram/sel_a[3] ), .Y(a[29]) );
  INVX1 \myram/m3/ta/t28/U1  ( .A(\myram/m3/dout[28] ), .Y(n435) );
  TBUFX2 \myram/m3/ta/t28/b1  ( .A(n435), .EN(\myram/sel_a[3] ), .Y(a[28]) );
  INVX1 \myram/m3/ta/t27/U1  ( .A(\myram/m3/dout[27] ), .Y(n434) );
  TBUFX2 \myram/m3/ta/t27/b1  ( .A(n434), .EN(\myram/sel_a[3] ), .Y(a[27]) );
  INVX1 \myram/m3/ta/t26/U1  ( .A(\myram/m3/dout[26] ), .Y(n433) );
  TBUFX2 \myram/m3/ta/t26/b1  ( .A(n433), .EN(\myram/sel_a[3] ), .Y(a[26]) );
  INVX1 \myram/m3/ta/t25/U1  ( .A(\myram/m3/dout[25] ), .Y(n432) );
  TBUFX2 \myram/m3/ta/t25/b1  ( .A(n432), .EN(\myram/sel_a[3] ), .Y(a[25]) );
  INVX1 \myram/m3/ta/t24/U1  ( .A(\myram/m3/dout[24] ), .Y(n431) );
  TBUFX2 \myram/m3/ta/t24/b1  ( .A(n431), .EN(\myram/sel_a[3] ), .Y(a[24]) );
  INVX1 \myram/m3/ta/t23/U1  ( .A(\myram/m3/dout[23] ), .Y(n430) );
  TBUFX2 \myram/m3/ta/t23/b1  ( .A(n430), .EN(\myram/sel_a[3] ), .Y(a[23]) );
  INVX1 \myram/m3/ta/t22/U1  ( .A(\myram/m3/dout[22] ), .Y(n429) );
  TBUFX2 \myram/m3/ta/t22/b1  ( .A(n429), .EN(\myram/sel_a[3] ), .Y(a[22]) );
  INVX1 \myram/m3/ta/t21/U1  ( .A(\myram/m3/dout[21] ), .Y(n428) );
  TBUFX2 \myram/m3/ta/t21/b1  ( .A(n428), .EN(\myram/sel_a[3] ), .Y(a[21]) );
  INVX1 \myram/m3/ta/t20/U1  ( .A(\myram/m3/dout[20] ), .Y(n427) );
  TBUFX2 \myram/m3/ta/t20/b1  ( .A(n427), .EN(\myram/sel_a[3] ), .Y(a[20]) );
  INVX1 \myram/m3/ta/t19/U1  ( .A(\myram/m3/dout[19] ), .Y(n426) );
  TBUFX2 \myram/m3/ta/t19/b1  ( .A(n426), .EN(\myram/sel_a[3] ), .Y(a[19]) );
  INVX1 \myram/m3/ta/t18/U1  ( .A(\myram/m3/dout[18] ), .Y(n425) );
  TBUFX2 \myram/m3/ta/t18/b1  ( .A(n425), .EN(\myram/sel_a[3] ), .Y(a[18]) );
  INVX1 \myram/m3/ta/t17/U1  ( .A(\myram/m3/dout[17] ), .Y(n424) );
  TBUFX2 \myram/m3/ta/t17/b1  ( .A(n424), .EN(\myram/sel_a[3] ), .Y(a[17]) );
  INVX1 \myram/m3/ta/t16/U1  ( .A(\myram/m3/dout[16] ), .Y(n423) );
  TBUFX2 \myram/m3/ta/t16/b1  ( .A(n423), .EN(\myram/sel_a[3] ), .Y(a[16]) );
  INVX1 \myram/m3/ta/t15/U1  ( .A(\myram/m3/dout[15] ), .Y(n422) );
  TBUFX2 \myram/m3/ta/t15/b1  ( .A(n422), .EN(\myram/sel_a[3] ), .Y(a[15]) );
  INVX1 \myram/m3/ta/t14/U1  ( .A(\myram/m3/dout[14] ), .Y(n421) );
  TBUFX2 \myram/m3/ta/t14/b1  ( .A(n421), .EN(\myram/sel_a[3] ), .Y(a[14]) );
  INVX1 \myram/m3/ta/t13/U1  ( .A(\myram/m3/dout[13] ), .Y(n420) );
  TBUFX2 \myram/m3/ta/t13/b1  ( .A(n420), .EN(n236), .Y(a[13]) );
  INVX1 \myram/m3/ta/t12/U1  ( .A(\myram/m3/dout[12] ), .Y(n419) );
  TBUFX2 \myram/m3/ta/t12/b1  ( .A(n419), .EN(n236), .Y(a[12]) );
  INVX1 \myram/m3/ta/t11/U1  ( .A(\myram/m3/dout[11] ), .Y(n418) );
  TBUFX2 \myram/m3/ta/t11/b1  ( .A(n418), .EN(n236), .Y(a[11]) );
  INVX1 \myram/m3/ta/t10/U1  ( .A(\myram/m3/dout[10] ), .Y(n417) );
  TBUFX2 \myram/m3/ta/t10/b1  ( .A(n417), .EN(n236), .Y(a[10]) );
  INVX1 \myram/m3/ta/t9/U1  ( .A(\myram/m3/dout[9] ), .Y(n416) );
  TBUFX2 \myram/m3/ta/t9/b1  ( .A(n416), .EN(n236), .Y(a[9]) );
  INVX1 \myram/m3/ta/t8/U1  ( .A(\myram/m3/dout[8] ), .Y(n415) );
  TBUFX2 \myram/m3/ta/t8/b1  ( .A(n415), .EN(n236), .Y(a[8]) );
  INVX1 \myram/m3/ta/t7/U1  ( .A(\myram/m3/dout[7] ), .Y(n414) );
  TBUFX2 \myram/m3/ta/t7/b1  ( .A(n414), .EN(n236), .Y(a[7]) );
  INVX1 \myram/m3/ta/t6/U1  ( .A(\myram/m3/dout[6] ), .Y(n413) );
  TBUFX2 \myram/m3/ta/t6/b1  ( .A(n413), .EN(n236), .Y(a[6]) );
  INVX1 \myram/m3/ta/t5/U1  ( .A(\myram/m3/dout[5] ), .Y(n412) );
  TBUFX2 \myram/m3/ta/t5/b1  ( .A(n412), .EN(n236), .Y(a[5]) );
  TBUFX2 \myram/m3/ta/t4/b1  ( .A(n443), .EN(n236), .Y(a[4]) );
  TBUFX2 \myram/m3/ta/t3/b1  ( .A(n442), .EN(n236), .Y(a[3]) );
  TBUFX2 \myram/m3/ta/t2/b1  ( .A(n441), .EN(n236), .Y(a[2]) );
  TBUFX2 \myram/m3/ta/t1/b1  ( .A(n440), .EN(n236), .Y(a[1]) );
  TBUFX2 \myram/m3/ta/t0/b1  ( .A(n439), .EN(n236), .Y(a[0]) );
  TBUFX2 \myram/m2/tb/t31/b1  ( .A(n406), .EN(n284), .Y(b[31]) );
  TBUFX2 \myram/m2/tb/t30/b1  ( .A(n405), .EN(n284), .Y(b[30]) );
  TBUFX2 \myram/m2/tb/t29/b1  ( .A(n404), .EN(n284), .Y(b[29]) );
  TBUFX2 \myram/m2/tb/t28/b1  ( .A(n403), .EN(n284), .Y(b[28]) );
  TBUFX2 \myram/m2/tb/t27/b1  ( .A(n402), .EN(n284), .Y(b[27]) );
  TBUFX2 \myram/m2/tb/t26/b1  ( .A(n401), .EN(n284), .Y(b[26]) );
  TBUFX2 \myram/m2/tb/t25/b1  ( .A(n400), .EN(n284), .Y(b[25]) );
  TBUFX2 \myram/m2/tb/t24/b1  ( .A(n399), .EN(n284), .Y(b[24]) );
  TBUFX2 \myram/m2/tb/t23/b1  ( .A(n398), .EN(n284), .Y(b[23]) );
  TBUFX2 \myram/m2/tb/t22/b1  ( .A(n397), .EN(n284), .Y(b[22]) );
  TBUFX2 \myram/m2/tb/t21/b1  ( .A(n396), .EN(n284), .Y(b[21]) );
  TBUFX2 \myram/m2/tb/t20/b1  ( .A(n395), .EN(n284), .Y(b[20]) );
  TBUFX2 \myram/m2/tb/t19/b1  ( .A(n394), .EN(n284), .Y(b[19]) );
  TBUFX2 \myram/m2/tb/t18/b1  ( .A(n393), .EN(n284), .Y(b[18]) );
  TBUFX2 \myram/m2/tb/t17/b1  ( .A(n392), .EN(n284), .Y(b[17]) );
  TBUFX2 \myram/m2/tb/t16/b1  ( .A(n391), .EN(n284), .Y(b[16]) );
  TBUFX2 \myram/m2/tb/t15/b1  ( .A(n390), .EN(n284), .Y(b[15]) );
  TBUFX2 \myram/m2/tb/t14/b1  ( .A(n389), .EN(n284), .Y(b[14]) );
  TBUFX2 \myram/m2/tb/t13/b1  ( .A(n388), .EN(n284), .Y(b[13]) );
  TBUFX2 \myram/m2/tb/t12/b1  ( .A(n387), .EN(n283), .Y(b[12]) );
  TBUFX2 \myram/m2/tb/t11/b1  ( .A(n386), .EN(n283), .Y(b[11]) );
  TBUFX2 \myram/m2/tb/t10/b1  ( .A(n385), .EN(n283), .Y(b[10]) );
  TBUFX2 \myram/m2/tb/t9/b1  ( .A(n384), .EN(n283), .Y(b[9]) );
  TBUFX2 \myram/m2/tb/t8/b1  ( .A(n383), .EN(n283), .Y(b[8]) );
  TBUFX2 \myram/m2/tb/t7/b1  ( .A(n382), .EN(n283), .Y(b[7]) );
  TBUFX2 \myram/m2/tb/t6/b1  ( .A(n381), .EN(n283), .Y(b[6]) );
  TBUFX2 \myram/m2/tb/t5/b1  ( .A(n380), .EN(n283), .Y(b[5]) );
  INVX1 \myram/m2/tb/t4/U1  ( .A(\myram/m2/dout[4] ), .Y(n411) );
  TBUFX2 \myram/m2/tb/t4/b1  ( .A(n411), .EN(n283), .Y(b[4]) );
  INVX1 \myram/m2/tb/t3/U1  ( .A(\myram/m2/dout[3] ), .Y(n410) );
  TBUFX2 \myram/m2/tb/t3/b1  ( .A(n410), .EN(n283), .Y(b[3]) );
  INVX1 \myram/m2/tb/t2/U1  ( .A(\myram/m2/dout[2] ), .Y(n409) );
  TBUFX2 \myram/m2/tb/t2/b1  ( .A(n409), .EN(n283), .Y(b[2]) );
  INVX1 \myram/m2/tb/t1/U1  ( .A(\myram/m2/dout[1] ), .Y(n408) );
  TBUFX2 \myram/m2/tb/t1/b1  ( .A(n408), .EN(n283), .Y(b[1]) );
  INVX1 \myram/m2/tb/t0/U1  ( .A(\myram/m2/dout[0] ), .Y(n407) );
  TBUFX2 \myram/m2/tb/t0/b1  ( .A(n407), .EN(n283), .Y(b[0]) );
  INVX1 \myram/m2/ta/t31/U1  ( .A(\myram/m2/dout[31] ), .Y(n406) );
  TBUFX2 \myram/m2/ta/t31/b1  ( .A(n406), .EN(\myram/sel_a[2] ), .Y(a[31]) );
  INVX1 \myram/m2/ta/t30/U1  ( .A(\myram/m2/dout[30] ), .Y(n405) );
  TBUFX2 \myram/m2/ta/t30/b1  ( .A(n405), .EN(\myram/sel_a[2] ), .Y(a[30]) );
  INVX1 \myram/m2/ta/t29/U1  ( .A(\myram/m2/dout[29] ), .Y(n404) );
  TBUFX2 \myram/m2/ta/t29/b1  ( .A(n404), .EN(\myram/sel_a[2] ), .Y(a[29]) );
  INVX1 \myram/m2/ta/t28/U1  ( .A(\myram/m2/dout[28] ), .Y(n403) );
  TBUFX2 \myram/m2/ta/t28/b1  ( .A(n403), .EN(\myram/sel_a[2] ), .Y(a[28]) );
  INVX1 \myram/m2/ta/t27/U1  ( .A(\myram/m2/dout[27] ), .Y(n402) );
  TBUFX2 \myram/m2/ta/t27/b1  ( .A(n402), .EN(\myram/sel_a[2] ), .Y(a[27]) );
  INVX1 \myram/m2/ta/t26/U1  ( .A(\myram/m2/dout[26] ), .Y(n401) );
  TBUFX2 \myram/m2/ta/t26/b1  ( .A(n401), .EN(\myram/sel_a[2] ), .Y(a[26]) );
  INVX1 \myram/m2/ta/t25/U1  ( .A(\myram/m2/dout[25] ), .Y(n400) );
  TBUFX2 \myram/m2/ta/t25/b1  ( .A(n400), .EN(\myram/sel_a[2] ), .Y(a[25]) );
  INVX1 \myram/m2/ta/t24/U1  ( .A(\myram/m2/dout[24] ), .Y(n399) );
  TBUFX2 \myram/m2/ta/t24/b1  ( .A(n399), .EN(\myram/sel_a[2] ), .Y(a[24]) );
  INVX1 \myram/m2/ta/t23/U1  ( .A(\myram/m2/dout[23] ), .Y(n398) );
  TBUFX2 \myram/m2/ta/t23/b1  ( .A(n398), .EN(\myram/sel_a[2] ), .Y(a[23]) );
  INVX1 \myram/m2/ta/t22/U1  ( .A(\myram/m2/dout[22] ), .Y(n397) );
  TBUFX2 \myram/m2/ta/t22/b1  ( .A(n397), .EN(\myram/sel_a[2] ), .Y(a[22]) );
  INVX1 \myram/m2/ta/t21/U1  ( .A(\myram/m2/dout[21] ), .Y(n396) );
  TBUFX2 \myram/m2/ta/t21/b1  ( .A(n396), .EN(\myram/sel_a[2] ), .Y(a[21]) );
  INVX1 \myram/m2/ta/t20/U1  ( .A(\myram/m2/dout[20] ), .Y(n395) );
  TBUFX2 \myram/m2/ta/t20/b1  ( .A(n395), .EN(\myram/sel_a[2] ), .Y(a[20]) );
  INVX1 \myram/m2/ta/t19/U1  ( .A(\myram/m2/dout[19] ), .Y(n394) );
  TBUFX2 \myram/m2/ta/t19/b1  ( .A(n394), .EN(\myram/sel_a[2] ), .Y(a[19]) );
  INVX1 \myram/m2/ta/t18/U1  ( .A(\myram/m2/dout[18] ), .Y(n393) );
  TBUFX2 \myram/m2/ta/t18/b1  ( .A(n393), .EN(\myram/sel_a[2] ), .Y(a[18]) );
  INVX1 \myram/m2/ta/t17/U1  ( .A(\myram/m2/dout[17] ), .Y(n392) );
  TBUFX2 \myram/m2/ta/t17/b1  ( .A(n392), .EN(\myram/sel_a[2] ), .Y(a[17]) );
  INVX1 \myram/m2/ta/t16/U1  ( .A(\myram/m2/dout[16] ), .Y(n391) );
  TBUFX2 \myram/m2/ta/t16/b1  ( .A(n391), .EN(\myram/sel_a[2] ), .Y(a[16]) );
  INVX1 \myram/m2/ta/t15/U1  ( .A(\myram/m2/dout[15] ), .Y(n390) );
  TBUFX2 \myram/m2/ta/t15/b1  ( .A(n390), .EN(\myram/sel_a[2] ), .Y(a[15]) );
  INVX1 \myram/m2/ta/t14/U1  ( .A(\myram/m2/dout[14] ), .Y(n389) );
  TBUFX2 \myram/m2/ta/t14/b1  ( .A(n389), .EN(\myram/sel_a[2] ), .Y(a[14]) );
  INVX1 \myram/m2/ta/t13/U1  ( .A(\myram/m2/dout[13] ), .Y(n388) );
  TBUFX2 \myram/m2/ta/t13/b1  ( .A(n388), .EN(n238), .Y(a[13]) );
  INVX1 \myram/m2/ta/t12/U1  ( .A(\myram/m2/dout[12] ), .Y(n387) );
  TBUFX2 \myram/m2/ta/t12/b1  ( .A(n387), .EN(n238), .Y(a[12]) );
  INVX1 \myram/m2/ta/t11/U1  ( .A(\myram/m2/dout[11] ), .Y(n386) );
  TBUFX2 \myram/m2/ta/t11/b1  ( .A(n386), .EN(n238), .Y(a[11]) );
  INVX1 \myram/m2/ta/t10/U1  ( .A(\myram/m2/dout[10] ), .Y(n385) );
  TBUFX2 \myram/m2/ta/t10/b1  ( .A(n385), .EN(n238), .Y(a[10]) );
  INVX1 \myram/m2/ta/t9/U1  ( .A(\myram/m2/dout[9] ), .Y(n384) );
  TBUFX2 \myram/m2/ta/t9/b1  ( .A(n384), .EN(n238), .Y(a[9]) );
  INVX1 \myram/m2/ta/t8/U1  ( .A(\myram/m2/dout[8] ), .Y(n383) );
  TBUFX2 \myram/m2/ta/t8/b1  ( .A(n383), .EN(n238), .Y(a[8]) );
  INVX1 \myram/m2/ta/t7/U1  ( .A(\myram/m2/dout[7] ), .Y(n382) );
  TBUFX2 \myram/m2/ta/t7/b1  ( .A(n382), .EN(n238), .Y(a[7]) );
  INVX1 \myram/m2/ta/t6/U1  ( .A(\myram/m2/dout[6] ), .Y(n381) );
  TBUFX2 \myram/m2/ta/t6/b1  ( .A(n381), .EN(n238), .Y(a[6]) );
  INVX1 \myram/m2/ta/t5/U1  ( .A(\myram/m2/dout[5] ), .Y(n380) );
  TBUFX2 \myram/m2/ta/t5/b1  ( .A(n380), .EN(n238), .Y(a[5]) );
  TBUFX2 \myram/m2/ta/t4/b1  ( .A(n411), .EN(n238), .Y(a[4]) );
  TBUFX2 \myram/m2/ta/t3/b1  ( .A(n410), .EN(n238), .Y(a[3]) );
  TBUFX2 \myram/m2/ta/t2/b1  ( .A(n409), .EN(n238), .Y(a[2]) );
  TBUFX2 \myram/m2/ta/t1/b1  ( .A(n408), .EN(n238), .Y(a[1]) );
  TBUFX2 \myram/m2/ta/t0/b1  ( .A(n407), .EN(n238), .Y(a[0]) );
  TBUFX2 \myram/m1/tb/t31/b1  ( .A(n374), .EN(n287), .Y(b[31]) );
  TBUFX2 \myram/m1/tb/t30/b1  ( .A(n373), .EN(n287), .Y(b[30]) );
  TBUFX2 \myram/m1/tb/t29/b1  ( .A(n372), .EN(n287), .Y(b[29]) );
  TBUFX2 \myram/m1/tb/t28/b1  ( .A(n371), .EN(n287), .Y(b[28]) );
  TBUFX2 \myram/m1/tb/t27/b1  ( .A(n370), .EN(n287), .Y(b[27]) );
  TBUFX2 \myram/m1/tb/t26/b1  ( .A(n369), .EN(n287), .Y(b[26]) );
  TBUFX2 \myram/m1/tb/t25/b1  ( .A(n368), .EN(n287), .Y(b[25]) );
  TBUFX2 \myram/m1/tb/t24/b1  ( .A(n367), .EN(n287), .Y(b[24]) );
  TBUFX2 \myram/m1/tb/t23/b1  ( .A(n366), .EN(n287), .Y(b[23]) );
  TBUFX2 \myram/m1/tb/t22/b1  ( .A(n365), .EN(n287), .Y(b[22]) );
  TBUFX2 \myram/m1/tb/t21/b1  ( .A(n364), .EN(n287), .Y(b[21]) );
  TBUFX2 \myram/m1/tb/t20/b1  ( .A(n363), .EN(n287), .Y(b[20]) );
  TBUFX2 \myram/m1/tb/t19/b1  ( .A(n362), .EN(n287), .Y(b[19]) );
  TBUFX2 \myram/m1/tb/t18/b1  ( .A(n361), .EN(n287), .Y(b[18]) );
  TBUFX2 \myram/m1/tb/t17/b1  ( .A(n360), .EN(n287), .Y(b[17]) );
  TBUFX2 \myram/m1/tb/t16/b1  ( .A(n359), .EN(n287), .Y(b[16]) );
  TBUFX2 \myram/m1/tb/t15/b1  ( .A(n358), .EN(n287), .Y(b[15]) );
  TBUFX2 \myram/m1/tb/t14/b1  ( .A(n357), .EN(n287), .Y(b[14]) );
  TBUFX2 \myram/m1/tb/t13/b1  ( .A(n356), .EN(n287), .Y(b[13]) );
  TBUFX2 \myram/m1/tb/t12/b1  ( .A(n355), .EN(n286), .Y(b[12]) );
  TBUFX2 \myram/m1/tb/t11/b1  ( .A(n354), .EN(n286), .Y(b[11]) );
  TBUFX2 \myram/m1/tb/t10/b1  ( .A(n353), .EN(n286), .Y(b[10]) );
  TBUFX2 \myram/m1/tb/t9/b1  ( .A(n352), .EN(n286), .Y(b[9]) );
  TBUFX2 \myram/m1/tb/t8/b1  ( .A(n351), .EN(n286), .Y(b[8]) );
  TBUFX2 \myram/m1/tb/t7/b1  ( .A(n350), .EN(n286), .Y(b[7]) );
  TBUFX2 \myram/m1/tb/t6/b1  ( .A(n349), .EN(n286), .Y(b[6]) );
  TBUFX2 \myram/m1/tb/t5/b1  ( .A(n348), .EN(n286), .Y(b[5]) );
  INVX1 \myram/m1/tb/t4/U1  ( .A(\myram/m1/dout[4] ), .Y(n379) );
  TBUFX2 \myram/m1/tb/t4/b1  ( .A(n379), .EN(n286), .Y(b[4]) );
  INVX1 \myram/m1/tb/t3/U1  ( .A(\myram/m1/dout[3] ), .Y(n378) );
  TBUFX2 \myram/m1/tb/t3/b1  ( .A(n378), .EN(n286), .Y(b[3]) );
  INVX1 \myram/m1/tb/t2/U1  ( .A(\myram/m1/dout[2] ), .Y(n377) );
  TBUFX2 \myram/m1/tb/t2/b1  ( .A(n377), .EN(n286), .Y(b[2]) );
  INVX1 \myram/m1/tb/t1/U1  ( .A(\myram/m1/dout[1] ), .Y(n376) );
  TBUFX2 \myram/m1/tb/t1/b1  ( .A(n376), .EN(n286), .Y(b[1]) );
  INVX1 \myram/m1/tb/t0/U1  ( .A(\myram/m1/dout[0] ), .Y(n375) );
  TBUFX2 \myram/m1/tb/t0/b1  ( .A(n375), .EN(n286), .Y(b[0]) );
  INVX1 \myram/m1/ta/t31/U1  ( .A(\myram/m1/dout[31] ), .Y(n374) );
  TBUFX2 \myram/m1/ta/t31/b1  ( .A(n374), .EN(\myram/sel_a[1] ), .Y(a[31]) );
  INVX1 \myram/m1/ta/t30/U1  ( .A(\myram/m1/dout[30] ), .Y(n373) );
  TBUFX2 \myram/m1/ta/t30/b1  ( .A(n373), .EN(\myram/sel_a[1] ), .Y(a[30]) );
  INVX1 \myram/m1/ta/t29/U1  ( .A(\myram/m1/dout[29] ), .Y(n372) );
  TBUFX2 \myram/m1/ta/t29/b1  ( .A(n372), .EN(\myram/sel_a[1] ), .Y(a[29]) );
  INVX1 \myram/m1/ta/t28/U1  ( .A(\myram/m1/dout[28] ), .Y(n371) );
  TBUFX2 \myram/m1/ta/t28/b1  ( .A(n371), .EN(\myram/sel_a[1] ), .Y(a[28]) );
  INVX1 \myram/m1/ta/t27/U1  ( .A(\myram/m1/dout[27] ), .Y(n370) );
  TBUFX2 \myram/m1/ta/t27/b1  ( .A(n370), .EN(\myram/sel_a[1] ), .Y(a[27]) );
  INVX1 \myram/m1/ta/t26/U1  ( .A(\myram/m1/dout[26] ), .Y(n369) );
  TBUFX2 \myram/m1/ta/t26/b1  ( .A(n369), .EN(\myram/sel_a[1] ), .Y(a[26]) );
  INVX1 \myram/m1/ta/t25/U1  ( .A(\myram/m1/dout[25] ), .Y(n368) );
  TBUFX2 \myram/m1/ta/t25/b1  ( .A(n368), .EN(\myram/sel_a[1] ), .Y(a[25]) );
  INVX1 \myram/m1/ta/t24/U1  ( .A(\myram/m1/dout[24] ), .Y(n367) );
  TBUFX2 \myram/m1/ta/t24/b1  ( .A(n367), .EN(\myram/sel_a[1] ), .Y(a[24]) );
  INVX1 \myram/m1/ta/t23/U1  ( .A(\myram/m1/dout[23] ), .Y(n366) );
  TBUFX2 \myram/m1/ta/t23/b1  ( .A(n366), .EN(\myram/sel_a[1] ), .Y(a[23]) );
  INVX1 \myram/m1/ta/t22/U1  ( .A(\myram/m1/dout[22] ), .Y(n365) );
  TBUFX2 \myram/m1/ta/t22/b1  ( .A(n365), .EN(\myram/sel_a[1] ), .Y(a[22]) );
  INVX1 \myram/m1/ta/t21/U1  ( .A(\myram/m1/dout[21] ), .Y(n364) );
  TBUFX2 \myram/m1/ta/t21/b1  ( .A(n364), .EN(\myram/sel_a[1] ), .Y(a[21]) );
  INVX1 \myram/m1/ta/t20/U1  ( .A(\myram/m1/dout[20] ), .Y(n363) );
  TBUFX2 \myram/m1/ta/t20/b1  ( .A(n363), .EN(\myram/sel_a[1] ), .Y(a[20]) );
  INVX1 \myram/m1/ta/t19/U1  ( .A(\myram/m1/dout[19] ), .Y(n362) );
  TBUFX2 \myram/m1/ta/t19/b1  ( .A(n362), .EN(\myram/sel_a[1] ), .Y(a[19]) );
  INVX1 \myram/m1/ta/t18/U1  ( .A(\myram/m1/dout[18] ), .Y(n361) );
  TBUFX2 \myram/m1/ta/t18/b1  ( .A(n361), .EN(\myram/sel_a[1] ), .Y(a[18]) );
  INVX1 \myram/m1/ta/t17/U1  ( .A(\myram/m1/dout[17] ), .Y(n360) );
  TBUFX2 \myram/m1/ta/t17/b1  ( .A(n360), .EN(\myram/sel_a[1] ), .Y(a[17]) );
  INVX1 \myram/m1/ta/t16/U1  ( .A(\myram/m1/dout[16] ), .Y(n359) );
  TBUFX2 \myram/m1/ta/t16/b1  ( .A(n359), .EN(\myram/sel_a[1] ), .Y(a[16]) );
  INVX1 \myram/m1/ta/t15/U1  ( .A(\myram/m1/dout[15] ), .Y(n358) );
  TBUFX2 \myram/m1/ta/t15/b1  ( .A(n358), .EN(\myram/sel_a[1] ), .Y(a[15]) );
  INVX1 \myram/m1/ta/t14/U1  ( .A(\myram/m1/dout[14] ), .Y(n357) );
  TBUFX2 \myram/m1/ta/t14/b1  ( .A(n357), .EN(\myram/sel_a[1] ), .Y(a[14]) );
  INVX1 \myram/m1/ta/t13/U1  ( .A(\myram/m1/dout[13] ), .Y(n356) );
  TBUFX2 \myram/m1/ta/t13/b1  ( .A(n356), .EN(n240), .Y(a[13]) );
  INVX1 \myram/m1/ta/t12/U1  ( .A(\myram/m1/dout[12] ), .Y(n355) );
  TBUFX2 \myram/m1/ta/t12/b1  ( .A(n355), .EN(n240), .Y(a[12]) );
  INVX1 \myram/m1/ta/t11/U1  ( .A(\myram/m1/dout[11] ), .Y(n354) );
  TBUFX2 \myram/m1/ta/t11/b1  ( .A(n354), .EN(n240), .Y(a[11]) );
  INVX1 \myram/m1/ta/t10/U1  ( .A(\myram/m1/dout[10] ), .Y(n353) );
  TBUFX2 \myram/m1/ta/t10/b1  ( .A(n353), .EN(n240), .Y(a[10]) );
  INVX1 \myram/m1/ta/t9/U1  ( .A(\myram/m1/dout[9] ), .Y(n352) );
  TBUFX2 \myram/m1/ta/t9/b1  ( .A(n352), .EN(n240), .Y(a[9]) );
  INVX1 \myram/m1/ta/t8/U1  ( .A(\myram/m1/dout[8] ), .Y(n351) );
  TBUFX2 \myram/m1/ta/t8/b1  ( .A(n351), .EN(n240), .Y(a[8]) );
  INVX1 \myram/m1/ta/t7/U1  ( .A(\myram/m1/dout[7] ), .Y(n350) );
  TBUFX2 \myram/m1/ta/t7/b1  ( .A(n350), .EN(n240), .Y(a[7]) );
  INVX1 \myram/m1/ta/t6/U1  ( .A(\myram/m1/dout[6] ), .Y(n349) );
  TBUFX2 \myram/m1/ta/t6/b1  ( .A(n349), .EN(n240), .Y(a[6]) );
  INVX1 \myram/m1/ta/t5/U1  ( .A(\myram/m1/dout[5] ), .Y(n348) );
  TBUFX2 \myram/m1/ta/t5/b1  ( .A(n348), .EN(n240), .Y(a[5]) );
  TBUFX2 \myram/m1/ta/t4/b1  ( .A(n379), .EN(n240), .Y(a[4]) );
  TBUFX2 \myram/m1/ta/t3/b1  ( .A(n378), .EN(n240), .Y(a[3]) );
  TBUFX2 \myram/m1/ta/t2/b1  ( .A(n377), .EN(n240), .Y(a[2]) );
  TBUFX2 \myram/m1/ta/t1/b1  ( .A(n376), .EN(n240), .Y(a[1]) );
  TBUFX2 \myram/m1/ta/t0/b1  ( .A(n375), .EN(n240), .Y(a[0]) );
  TBUFX2 \myram/m0/tb/t31/b1  ( .A(n342), .EN(n290), .Y(b[31]) );
  TBUFX2 \myram/m0/tb/t30/b1  ( .A(n341), .EN(n290), .Y(b[30]) );
  TBUFX2 \myram/m0/tb/t29/b1  ( .A(n340), .EN(n290), .Y(b[29]) );
  TBUFX2 \myram/m0/tb/t28/b1  ( .A(n339), .EN(n290), .Y(b[28]) );
  TBUFX2 \myram/m0/tb/t27/b1  ( .A(n338), .EN(n290), .Y(b[27]) );
  TBUFX2 \myram/m0/tb/t26/b1  ( .A(n337), .EN(n290), .Y(b[26]) );
  TBUFX2 \myram/m0/tb/t25/b1  ( .A(n336), .EN(n290), .Y(b[25]) );
  TBUFX2 \myram/m0/tb/t24/b1  ( .A(n335), .EN(n290), .Y(b[24]) );
  TBUFX2 \myram/m0/tb/t23/b1  ( .A(n334), .EN(n290), .Y(b[23]) );
  TBUFX2 \myram/m0/tb/t22/b1  ( .A(n333), .EN(n290), .Y(b[22]) );
  TBUFX2 \myram/m0/tb/t21/b1  ( .A(n332), .EN(n290), .Y(b[21]) );
  TBUFX2 \myram/m0/tb/t20/b1  ( .A(n331), .EN(n290), .Y(b[20]) );
  TBUFX2 \myram/m0/tb/t19/b1  ( .A(n330), .EN(n290), .Y(b[19]) );
  TBUFX2 \myram/m0/tb/t18/b1  ( .A(n329), .EN(n290), .Y(b[18]) );
  TBUFX2 \myram/m0/tb/t17/b1  ( .A(n328), .EN(n290), .Y(b[17]) );
  TBUFX2 \myram/m0/tb/t16/b1  ( .A(n327), .EN(n290), .Y(b[16]) );
  TBUFX2 \myram/m0/tb/t15/b1  ( .A(n326), .EN(n290), .Y(b[15]) );
  TBUFX2 \myram/m0/tb/t14/b1  ( .A(n325), .EN(n290), .Y(b[14]) );
  TBUFX2 \myram/m0/tb/t13/b1  ( .A(n324), .EN(n290), .Y(b[13]) );
  TBUFX2 \myram/m0/tb/t12/b1  ( .A(n323), .EN(n289), .Y(b[12]) );
  TBUFX2 \myram/m0/tb/t11/b1  ( .A(n322), .EN(n289), .Y(b[11]) );
  TBUFX2 \myram/m0/tb/t10/b1  ( .A(n321), .EN(n289), .Y(b[10]) );
  TBUFX2 \myram/m0/tb/t9/b1  ( .A(n320), .EN(n289), .Y(b[9]) );
  TBUFX2 \myram/m0/tb/t8/b1  ( .A(n319), .EN(n289), .Y(b[8]) );
  TBUFX2 \myram/m0/tb/t7/b1  ( .A(n318), .EN(n289), .Y(b[7]) );
  TBUFX2 \myram/m0/tb/t6/b1  ( .A(n317), .EN(n289), .Y(b[6]) );
  TBUFX2 \myram/m0/tb/t5/b1  ( .A(n316), .EN(n289), .Y(b[5]) );
  INVX1 \myram/m0/tb/t4/U1  ( .A(\myram/m0/dout[4] ), .Y(n347) );
  TBUFX2 \myram/m0/tb/t4/b1  ( .A(n347), .EN(n289), .Y(b[4]) );
  INVX1 \myram/m0/tb/t3/U1  ( .A(\myram/m0/dout[3] ), .Y(n346) );
  TBUFX2 \myram/m0/tb/t3/b1  ( .A(n346), .EN(n289), .Y(b[3]) );
  INVX1 \myram/m0/tb/t2/U1  ( .A(\myram/m0/dout[2] ), .Y(n345) );
  TBUFX2 \myram/m0/tb/t2/b1  ( .A(n345), .EN(n289), .Y(b[2]) );
  INVX1 \myram/m0/tb/t1/U1  ( .A(\myram/m0/dout[1] ), .Y(n344) );
  TBUFX2 \myram/m0/tb/t1/b1  ( .A(n344), .EN(n289), .Y(b[1]) );
  INVX1 \myram/m0/tb/t0/U1  ( .A(\myram/m0/dout[0] ), .Y(n343) );
  TBUFX2 \myram/m0/tb/t0/b1  ( .A(n343), .EN(n289), .Y(b[0]) );
  INVX1 \myram/m0/ta/t31/U1  ( .A(\myram/m0/dout[31] ), .Y(n342) );
  TBUFX2 \myram/m0/ta/t31/b1  ( .A(n342), .EN(\myram/sel_a[0] ), .Y(a[31]) );
  INVX1 \myram/m0/ta/t30/U1  ( .A(\myram/m0/dout[30] ), .Y(n341) );
  TBUFX2 \myram/m0/ta/t30/b1  ( .A(n341), .EN(\myram/sel_a[0] ), .Y(a[30]) );
  INVX1 \myram/m0/ta/t29/U1  ( .A(\myram/m0/dout[29] ), .Y(n340) );
  TBUFX2 \myram/m0/ta/t29/b1  ( .A(n340), .EN(\myram/sel_a[0] ), .Y(a[29]) );
  INVX1 \myram/m0/ta/t28/U1  ( .A(\myram/m0/dout[28] ), .Y(n339) );
  TBUFX2 \myram/m0/ta/t28/b1  ( .A(n339), .EN(\myram/sel_a[0] ), .Y(a[28]) );
  INVX1 \myram/m0/ta/t27/U1  ( .A(\myram/m0/dout[27] ), .Y(n338) );
  TBUFX2 \myram/m0/ta/t27/b1  ( .A(n338), .EN(\myram/sel_a[0] ), .Y(a[27]) );
  INVX1 \myram/m0/ta/t26/U1  ( .A(\myram/m0/dout[26] ), .Y(n337) );
  TBUFX2 \myram/m0/ta/t26/b1  ( .A(n337), .EN(\myram/sel_a[0] ), .Y(a[26]) );
  INVX1 \myram/m0/ta/t25/U1  ( .A(\myram/m0/dout[25] ), .Y(n336) );
  TBUFX2 \myram/m0/ta/t25/b1  ( .A(n336), .EN(\myram/sel_a[0] ), .Y(a[25]) );
  INVX1 \myram/m0/ta/t24/U1  ( .A(\myram/m0/dout[24] ), .Y(n335) );
  TBUFX2 \myram/m0/ta/t24/b1  ( .A(n335), .EN(\myram/sel_a[0] ), .Y(a[24]) );
  INVX1 \myram/m0/ta/t23/U1  ( .A(\myram/m0/dout[23] ), .Y(n334) );
  TBUFX2 \myram/m0/ta/t23/b1  ( .A(n334), .EN(\myram/sel_a[0] ), .Y(a[23]) );
  INVX1 \myram/m0/ta/t22/U1  ( .A(\myram/m0/dout[22] ), .Y(n333) );
  TBUFX2 \myram/m0/ta/t22/b1  ( .A(n333), .EN(\myram/sel_a[0] ), .Y(a[22]) );
  INVX1 \myram/m0/ta/t21/U1  ( .A(\myram/m0/dout[21] ), .Y(n332) );
  TBUFX2 \myram/m0/ta/t21/b1  ( .A(n332), .EN(\myram/sel_a[0] ), .Y(a[21]) );
  INVX1 \myram/m0/ta/t20/U1  ( .A(\myram/m0/dout[20] ), .Y(n331) );
  TBUFX2 \myram/m0/ta/t20/b1  ( .A(n331), .EN(\myram/sel_a[0] ), .Y(a[20]) );
  INVX1 \myram/m0/ta/t19/U1  ( .A(\myram/m0/dout[19] ), .Y(n330) );
  TBUFX2 \myram/m0/ta/t19/b1  ( .A(n330), .EN(\myram/sel_a[0] ), .Y(a[19]) );
  INVX1 \myram/m0/ta/t18/U1  ( .A(\myram/m0/dout[18] ), .Y(n329) );
  TBUFX2 \myram/m0/ta/t18/b1  ( .A(n329), .EN(\myram/sel_a[0] ), .Y(a[18]) );
  INVX1 \myram/m0/ta/t17/U1  ( .A(\myram/m0/dout[17] ), .Y(n328) );
  TBUFX2 \myram/m0/ta/t17/b1  ( .A(n328), .EN(\myram/sel_a[0] ), .Y(a[17]) );
  INVX1 \myram/m0/ta/t16/U1  ( .A(\myram/m0/dout[16] ), .Y(n327) );
  TBUFX2 \myram/m0/ta/t16/b1  ( .A(n327), .EN(\myram/sel_a[0] ), .Y(a[16]) );
  INVX1 \myram/m0/ta/t15/U1  ( .A(\myram/m0/dout[15] ), .Y(n326) );
  TBUFX2 \myram/m0/ta/t15/b1  ( .A(n326), .EN(n242), .Y(a[15]) );
  INVX1 \myram/m0/ta/t14/U1  ( .A(\myram/m0/dout[14] ), .Y(n325) );
  TBUFX2 \myram/m0/ta/t14/b1  ( .A(n325), .EN(\myram/sel_a[0] ), .Y(a[14]) );
  INVX1 \myram/m0/ta/t13/U1  ( .A(\myram/m0/dout[13] ), .Y(n324) );
  TBUFX2 \myram/m0/ta/t13/b1  ( .A(n324), .EN(n242), .Y(a[13]) );
  INVX1 \myram/m0/ta/t12/U1  ( .A(\myram/m0/dout[12] ), .Y(n323) );
  TBUFX2 \myram/m0/ta/t12/b1  ( .A(n323), .EN(n242), .Y(a[12]) );
  INVX1 \myram/m0/ta/t11/U1  ( .A(\myram/m0/dout[11] ), .Y(n322) );
  TBUFX2 \myram/m0/ta/t11/b1  ( .A(n322), .EN(n242), .Y(a[11]) );
  INVX1 \myram/m0/ta/t10/U1  ( .A(\myram/m0/dout[10] ), .Y(n321) );
  TBUFX2 \myram/m0/ta/t10/b1  ( .A(n321), .EN(n242), .Y(a[10]) );
  INVX1 \myram/m0/ta/t9/U1  ( .A(\myram/m0/dout[9] ), .Y(n320) );
  TBUFX2 \myram/m0/ta/t9/b1  ( .A(n320), .EN(n242), .Y(a[9]) );
  INVX1 \myram/m0/ta/t8/U1  ( .A(\myram/m0/dout[8] ), .Y(n319) );
  TBUFX2 \myram/m0/ta/t8/b1  ( .A(n319), .EN(n242), .Y(a[8]) );
  INVX1 \myram/m0/ta/t7/U1  ( .A(\myram/m0/dout[7] ), .Y(n318) );
  TBUFX2 \myram/m0/ta/t7/b1  ( .A(n318), .EN(n242), .Y(a[7]) );
  INVX1 \myram/m0/ta/t6/U1  ( .A(\myram/m0/dout[6] ), .Y(n317) );
  TBUFX2 \myram/m0/ta/t6/b1  ( .A(n317), .EN(n242), .Y(a[6]) );
  INVX1 \myram/m0/ta/t5/U1  ( .A(\myram/m0/dout[5] ), .Y(n316) );
  TBUFX2 \myram/m0/ta/t5/b1  ( .A(n316), .EN(n242), .Y(a[5]) );
  TBUFX2 \myram/m0/ta/t4/b1  ( .A(n347), .EN(n242), .Y(a[4]) );
  TBUFX2 \myram/m0/ta/t3/b1  ( .A(n346), .EN(n242), .Y(a[3]) );
  TBUFX2 \myram/m0/ta/t2/b1  ( .A(n345), .EN(n242), .Y(a[2]) );
  TBUFX2 \myram/m0/ta/t1/b1  ( .A(n344), .EN(n242), .Y(a[1]) );
  AND2X1 U26 ( .A(addr_s[3]), .B(write_en), .Y(\myram/ds/en1 ) );
  BUFX2 U27 ( .A(b[2]), .Y(n25) );
  AND2X1 U28 ( .A(addr_s[2]), .B(n110), .Y(\myram/ds/d0/en1 ) );
  INVX1 U29 ( .A(\myram/ds/en1 ), .Y(n841) );
  OR2X1 U30 ( .A(n104), .B(n105), .Y(n4) );
  BUFX4 U31 ( .A(b[1]), .Y(n62) );
  INVX1 U32 ( .A(\myram/db/en1 ), .Y(n840) );
  AND2X1 U33 ( .A(code[15]), .B(n125), .Y(n2169) );
  AND2X1 U34 ( .A(alu_s[9]), .B(n315), .Y(mem_s[9]) );
  BUFX2 U35 ( .A(n1001), .Y(n26) );
  INVX1 U36 ( .A(n26), .Y(\myalu/s10[0] ) );
  BUFX2 U37 ( .A(n1003), .Y(n27) );
  INVX1 U38 ( .A(n27), .Y(\myalu/s10[2] ) );
  BUFX2 U39 ( .A(n1004), .Y(n28) );
  INVX1 U40 ( .A(n28), .Y(\myalu/s10[3] ) );
  BUFX2 U41 ( .A(n1005), .Y(n29) );
  INVX1 U42 ( .A(n29), .Y(\myalu/s10[4] ) );
  BUFX2 U43 ( .A(n1006), .Y(n30) );
  INVX1 U44 ( .A(n30), .Y(\myalu/s10[5] ) );
  BUFX2 U45 ( .A(n1007), .Y(n31) );
  INVX1 U46 ( .A(n31), .Y(\myalu/s10[6] ) );
  BUFX2 U47 ( .A(n1008), .Y(n32) );
  INVX1 U48 ( .A(n32), .Y(\myalu/s10[7] ) );
  BUFX2 U49 ( .A(n1022), .Y(n33) );
  INVX1 U50 ( .A(n33), .Y(\myalu/s10[21] ) );
  BUFX2 U51 ( .A(n1023), .Y(n34) );
  INVX1 U52 ( .A(n34), .Y(\myalu/s10[22] ) );
  BUFX2 U53 ( .A(n1024), .Y(n35) );
  INVX1 U54 ( .A(n35), .Y(\myalu/s10[23] ) );
  BUFX2 U55 ( .A(n1026), .Y(n36) );
  INVX1 U56 ( .A(n36), .Y(\myalu/s10[25] ) );
  BUFX2 U57 ( .A(n1029), .Y(n37) );
  INVX1 U58 ( .A(n37), .Y(\myalu/s10[28] ) );
  BUFX2 U59 ( .A(n1030), .Y(n38) );
  INVX1 U60 ( .A(n38), .Y(\myalu/s10[29] ) );
  BUFX2 U61 ( .A(n1073), .Y(n39) );
  INVX1 U62 ( .A(n39), .Y(alu_s[8]) );
  BUFX2 U63 ( .A(n1075), .Y(n40) );
  INVX1 U64 ( .A(n40), .Y(alu_s[10]) );
  BUFX2 U65 ( .A(n1076), .Y(n41) );
  INVX1 U66 ( .A(n41), .Y(alu_s[11]) );
  BUFX2 U67 ( .A(n1077), .Y(n42) );
  INVX1 U68 ( .A(n42), .Y(alu_s[12]) );
  BUFX2 U69 ( .A(n1078), .Y(n43) );
  INVX1 U70 ( .A(n43), .Y(alu_s[13]) );
  BUFX2 U71 ( .A(n1079), .Y(n44) );
  INVX1 U72 ( .A(n44), .Y(alu_s[14]) );
  BUFX2 U73 ( .A(n1080), .Y(n45) );
  INVX1 U74 ( .A(n45), .Y(alu_s[15]) );
  BUFX2 U75 ( .A(n1081), .Y(n46) );
  INVX1 U76 ( .A(n46), .Y(alu_s[16]) );
  BUFX2 U77 ( .A(n1082), .Y(n47) );
  INVX1 U78 ( .A(n47), .Y(alu_s[17]) );
  BUFX2 U79 ( .A(n1083), .Y(n48) );
  INVX1 U80 ( .A(n48), .Y(alu_s[18]) );
  BUFX2 U81 ( .A(n1084), .Y(n49) );
  INVX1 U82 ( .A(n49), .Y(alu_s[19]) );
  BUFX2 U83 ( .A(n1085), .Y(n50) );
  INVX1 U84 ( .A(n50), .Y(alu_s[20]) );
  BUFX2 U85 ( .A(n1086), .Y(n51) );
  INVX1 U86 ( .A(n51), .Y(alu_s[21]) );
  BUFX2 U87 ( .A(n1087), .Y(n52) );
  INVX1 U88 ( .A(n52), .Y(alu_s[22]) );
  BUFX2 U89 ( .A(n1088), .Y(n53) );
  INVX1 U90 ( .A(n53), .Y(alu_s[23]) );
  BUFX2 U91 ( .A(n1089), .Y(n54) );
  INVX1 U92 ( .A(n54), .Y(alu_s[24]) );
  BUFX2 U93 ( .A(n1090), .Y(n55) );
  INVX1 U94 ( .A(n55), .Y(alu_s[25]) );
  BUFX2 U95 ( .A(n1091), .Y(n56) );
  INVX1 U96 ( .A(n56), .Y(alu_s[26]) );
  BUFX2 U97 ( .A(n1092), .Y(n57) );
  INVX1 U98 ( .A(n57), .Y(alu_s[27]) );
  BUFX2 U99 ( .A(n1093), .Y(n58) );
  INVX1 U100 ( .A(n58), .Y(alu_s[28]) );
  BUFX2 U101 ( .A(n1094), .Y(n59) );
  INVX1 U102 ( .A(n59), .Y(alu_s[29]) );
  BUFX2 U103 ( .A(n1095), .Y(n60) );
  INVX1 U104 ( .A(n60), .Y(alu_s[30]) );
  AND2X1 U105 ( .A(code[15]), .B(alu_op[1]), .Y(\myctl/n5 ) );
  INVX1 U106 ( .A(\myctl/n5 ), .Y(n61) );
  BUFX2 U107 ( .A(n1002), .Y(n63) );
  INVX1 U108 ( .A(n63), .Y(\myalu/s10[1] ) );
  BUFX2 U109 ( .A(n1021), .Y(n64) );
  INVX1 U110 ( .A(n64), .Y(\myalu/s10[20] ) );
  BUFX2 U111 ( .A(n960), .Y(n65) );
  INVX1 U112 ( .A(n65), .Y(\mypc/temp_pc1[0] ) );
  BUFX2 U113 ( .A(n1020), .Y(n66) );
  INVX1 U114 ( .A(n66), .Y(\myalu/s10[19] ) );
  BUFX2 U115 ( .A(n1017), .Y(n67) );
  INVX1 U116 ( .A(n67), .Y(\myalu/s10[16] ) );
  BUFX2 U117 ( .A(n968), .Y(n68) );
  INVX1 U118 ( .A(n68), .Y(\mypc/temp_pc1[7] ) );
  BUFX2 U119 ( .A(n1028), .Y(n69) );
  INVX1 U120 ( .A(n69), .Y(\myalu/s10[27] ) );
  BUFX2 U121 ( .A(n1016), .Y(n70) );
  INVX1 U122 ( .A(n70), .Y(\myalu/s10[15] ) );
  BUFX2 U123 ( .A(n967), .Y(n71) );
  INVX1 U124 ( .A(n71), .Y(\mypc/temp_pc1[6] ) );
  BUFX2 U125 ( .A(n1027), .Y(n72) );
  INVX1 U126 ( .A(n72), .Y(\myalu/s10[26] ) );
  BUFX2 U127 ( .A(n1015), .Y(n73) );
  INVX1 U128 ( .A(n73), .Y(\myalu/s10[14] ) );
  BUFX2 U129 ( .A(n966), .Y(n74) );
  INVX1 U130 ( .A(n74), .Y(\mypc/temp_pc1[5] ) );
  BUFX2 U131 ( .A(n1025), .Y(n75) );
  INVX1 U132 ( .A(n75), .Y(\myalu/s10[24] ) );
  BUFX2 U133 ( .A(n1014), .Y(n76) );
  INVX1 U134 ( .A(n76), .Y(\myalu/s10[13] ) );
  AND2X1 U135 ( .A(a[3]), .B(\myalu/myadder/xb[3] ), .Y(n859) );
  INVX1 U136 ( .A(n859), .Y(n77) );
  AND2X1 U137 ( .A(a[22]), .B(\myalu/myadder/xb[22] ), .Y(n916) );
  INVX1 U138 ( .A(n916), .Y(n78) );
  AND2X1 U139 ( .A(a[28]), .B(\myalu/myadder/xb[28] ), .Y(n934) );
  INVX1 U140 ( .A(n934), .Y(n79) );
  BUFX2 U141 ( .A(n965), .Y(n80) );
  INVX1 U142 ( .A(n80), .Y(\mypc/temp_pc1[4] ) );
  BUFX2 U143 ( .A(n1019), .Y(n81) );
  INVX1 U144 ( .A(n81), .Y(\myalu/s10[18] ) );
  BUFX2 U145 ( .A(n1013), .Y(n82) );
  INVX1 U146 ( .A(n82), .Y(\myalu/s10[12] ) );
  AND2X1 U147 ( .A(a[2]), .B(\myalu/myadder/xb[2] ), .Y(n856) );
  INVX1 U148 ( .A(n856), .Y(n83) );
  AND2X1 U149 ( .A(a[21]), .B(\myalu/myadder/xb[21] ), .Y(n913) );
  INVX1 U150 ( .A(n913), .Y(n84) );
  AND2X1 U151 ( .A(a[18]), .B(\myalu/myadder/xb[18] ), .Y(n904) );
  INVX1 U152 ( .A(n904), .Y(n85) );
  AND2X1 U153 ( .A(a[15]), .B(\myalu/myadder/xb[15] ), .Y(n895) );
  INVX1 U154 ( .A(n895), .Y(n86) );
  AND2X1 U155 ( .A(a[12]), .B(\myalu/myadder/xb[12] ), .Y(n886) );
  INVX1 U156 ( .A(n886), .Y(n87) );
  AND2X1 U157 ( .A(a[9]), .B(\myalu/myadder/xb[9] ), .Y(n877) );
  INVX1 U158 ( .A(n877), .Y(n88) );
  AND2X1 U159 ( .A(a[25]), .B(\myalu/myadder/xb[25] ), .Y(n925) );
  INVX1 U160 ( .A(n925), .Y(n89) );
  AND2X1 U161 ( .A(a[6]), .B(\myalu/myadder/xb[6] ), .Y(n868) );
  INVX1 U162 ( .A(n868), .Y(n90) );
  AND2X1 U163 ( .A(a[29]), .B(\myalu/myadder/xb[29] ), .Y(n937) );
  INVX1 U164 ( .A(n937), .Y(n91) );
  BUFX2 U165 ( .A(n964), .Y(n92) );
  INVX1 U166 ( .A(n92), .Y(\mypc/temp_pc1[3] ) );
  BUFX2 U167 ( .A(n1018), .Y(n93) );
  INVX1 U168 ( .A(n93), .Y(\myalu/s10[17] ) );
  BUFX2 U169 ( .A(n1012), .Y(n94) );
  INVX1 U170 ( .A(n94), .Y(\myalu/s10[11] ) );
  AND2X1 U171 ( .A(a[4]), .B(\myalu/myadder/xb[4] ), .Y(n862) );
  INVX1 U172 ( .A(n862), .Y(n95) );
  AND2X1 U173 ( .A(a[1]), .B(\myalu/myadder/xb[1] ), .Y(n853) );
  INVX1 U174 ( .A(n853), .Y(n96) );
  AND2X1 U175 ( .A(a[19]), .B(\myalu/myadder/xb[19] ), .Y(n907) );
  INVX1 U176 ( .A(n907), .Y(n97) );
  AND2X1 U177 ( .A(a[16]), .B(\myalu/myadder/xb[16] ), .Y(n898) );
  INVX1 U178 ( .A(n898), .Y(n98) );
  AND2X1 U179 ( .A(a[13]), .B(\myalu/myadder/xb[13] ), .Y(n889) );
  INVX1 U180 ( .A(n889), .Y(n99) );
  AND2X1 U181 ( .A(a[10]), .B(\myalu/myadder/xb[10] ), .Y(n880) );
  INVX1 U182 ( .A(n880), .Y(n100) );
  AND2X1 U183 ( .A(a[23]), .B(\myalu/myadder/xb[23] ), .Y(n919) );
  INVX1 U184 ( .A(n919), .Y(n101) );
  AND2X1 U185 ( .A(a[26]), .B(\myalu/myadder/xb[26] ), .Y(n928) );
  INVX1 U186 ( .A(n928), .Y(n102) );
  AND2X1 U187 ( .A(a[7]), .B(\myalu/myadder/xb[7] ), .Y(n871) );
  INVX1 U188 ( .A(n871), .Y(n103) );
  BUFX2 U189 ( .A(n5), .Y(n104) );
  BUFX2 U190 ( .A(n6), .Y(n105) );
  BUFX2 U191 ( .A(n963), .Y(n106) );
  INVX1 U192 ( .A(n106), .Y(\mypc/temp_pc1[2] ) );
  BUFX2 U193 ( .A(n1011), .Y(n107) );
  INVX1 U194 ( .A(n107), .Y(\myalu/s10[10] ) );
  BUFX2 U195 ( .A(n1031), .Y(n108) );
  INVX1 U196 ( .A(n108), .Y(\myalu/s10[30] ) );
  BUFX2 U197 ( .A(n1096), .Y(n109) );
  INVX1 U198 ( .A(n109), .Y(alu_s[31]) );
  OR2X1 U199 ( .A(addr_s[3]), .B(n2169), .Y(\myram/ds/en0 ) );
  INVX1 U200 ( .A(\myram/ds/en0 ), .Y(n110) );
  AND2X1 U201 ( .A(a[20]), .B(\myalu/myadder/xb[20] ), .Y(n910) );
  INVX1 U202 ( .A(n910), .Y(n111) );
  AND2X1 U203 ( .A(a[17]), .B(\myalu/myadder/xb[17] ), .Y(n901) );
  INVX1 U204 ( .A(n901), .Y(n112) );
  AND2X1 U205 ( .A(a[14]), .B(\myalu/myadder/xb[14] ), .Y(n892) );
  INVX1 U206 ( .A(n892), .Y(n113) );
  AND2X1 U207 ( .A(a[11]), .B(\myalu/myadder/xb[11] ), .Y(n883) );
  INVX1 U208 ( .A(n883), .Y(n114) );
  AND2X1 U209 ( .A(a[5]), .B(\myalu/myadder/xb[5] ), .Y(n865) );
  INVX1 U210 ( .A(n865), .Y(n115) );
  AND2X1 U211 ( .A(a[24]), .B(\myalu/myadder/xb[24] ), .Y(n922) );
  INVX1 U212 ( .A(n922), .Y(n116) );
  AND2X1 U213 ( .A(a[0]), .B(\myalu/myadder/xb[0] ), .Y(n850) );
  INVX1 U214 ( .A(n850), .Y(n117) );
  AND2X1 U215 ( .A(a[27]), .B(\myalu/myadder/xb[27] ), .Y(n931) );
  INVX1 U216 ( .A(n931), .Y(n118) );
  AND2X1 U217 ( .A(a[8]), .B(\myalu/myadder/xb[8] ), .Y(n874) );
  INVX1 U218 ( .A(n874), .Y(n119) );
  AND2X1 U219 ( .A(a[30]), .B(\myalu/myadder/xb[30] ), .Y(n940) );
  INVX1 U220 ( .A(n940), .Y(n120) );
  BUFX2 U221 ( .A(n962), .Y(n121) );
  INVX1 U222 ( .A(n121), .Y(\mypc/temp_pc1[1] ) );
  BUFX2 U223 ( .A(n1009), .Y(n122) );
  INVX1 U224 ( .A(n122), .Y(\myalu/s10[8] ) );
  BUFX2 U225 ( .A(n1032), .Y(n123) );
  INVX1 U226 ( .A(n123), .Y(\myalu/s10[31] ) );
  INVX1 U227 ( .A(n2169), .Y(write_en) );
  BUFX2 U228 ( .A(\myctl/n4 ), .Y(n125) );
  AND2X1 U229 ( .A(code[15]), .B(n314), .Y(\myctl/n6 ) );
  INVX1 U230 ( .A(\myctl/n6 ), .Y(n126) );
  AND2X1 U231 ( .A(alu_s[31]), .B(n315), .Y(mem_s[31]) );
  AND2X1 U232 ( .A(alu_s[31]), .B(n315), .Y(n132) );
  AND2X1 U233 ( .A(alu_s[31]), .B(n315), .Y(n128) );
  INVX1 U234 ( .A(n279), .Y(n277) );
  INVX1 U235 ( .A(n255), .Y(n253) );
  INVX1 U236 ( .A(n267), .Y(n265) );
  INVX1 U237 ( .A(n288), .Y(n286) );
  INVX1 U238 ( .A(n285), .Y(n283) );
  INVX1 U239 ( .A(n282), .Y(n280) );
  INVX1 U240 ( .A(n276), .Y(n274) );
  INVX1 U241 ( .A(n273), .Y(n271) );
  INVX1 U242 ( .A(n270), .Y(n268) );
  INVX1 U243 ( .A(n264), .Y(n262) );
  INVX1 U244 ( .A(n261), .Y(n259) );
  INVX1 U245 ( .A(n258), .Y(n256) );
  INVX1 U246 ( .A(n252), .Y(n250) );
  INVX1 U247 ( .A(n249), .Y(n247) );
  INVX1 U248 ( .A(n246), .Y(n244) );
  AND2X1 U249 ( .A(alu_s[30]), .B(n315), .Y(mem_s[30]) );
  BUFX2 U250 ( .A(addr_b[0]), .Y(n205) );
  BUFX2 U251 ( .A(addr_b[1]), .Y(n206) );
  INVX1 U252 ( .A(\myalu/myadder/myadder/c9 ), .Y(n875) );
  INVX1 U253 ( .A(\myalu/myadder/myadder/c5 ), .Y(n863) );
  INVX1 U254 ( .A(\myalu/myadder/myadder/c23 ), .Y(n917) );
  INVX1 U255 ( .A(\myalu/myadder/myadder/c12 ), .Y(n884) );
  INVX1 U256 ( .A(\myalu/myadder/myadder/c16 ), .Y(n896) );
  INVX1 U257 ( .A(\myalu/myadder/myadder/c20 ), .Y(n908) );
  INVX1 U258 ( .A(\myalu/myadder/myadder/c3 ), .Y(n857) );
  INVX1 U259 ( .A(\myalu/myadder/myadder/c6 ), .Y(n866) );
  INVX1 U260 ( .A(\myalu/myadder/myadder/c24 ), .Y(n920) );
  INVX1 U261 ( .A(\myalu/myadder/myadder/c10 ), .Y(n878) );
  INVX1 U262 ( .A(\myalu/myadder/myadder/c13 ), .Y(n887) );
  INVX1 U263 ( .A(\myalu/myadder/myadder/c17 ), .Y(n899) );
  INVX1 U264 ( .A(\myalu/myadder/myadder/c2 ), .Y(n854) );
  INVX1 U265 ( .A(\myalu/myadder/myadder/c26 ), .Y(n926) );
  INVX1 U266 ( .A(\myalu/myadder/myadder/c22 ), .Y(n914) );
  INVX1 U267 ( .A(\myalu/myadder/myadder/c11 ), .Y(n881) );
  INVX1 U268 ( .A(\myalu/myadder/myadder/c15 ), .Y(n893) );
  INVX1 U269 ( .A(\myalu/myadder/myadder/c19 ), .Y(n905) );
  INVX1 U270 ( .A(\myalu/myadder/myadder/c4 ), .Y(n860) );
  INVX1 U271 ( .A(\myalu/myadder/myadder/c7 ), .Y(n869) );
  INVX1 U272 ( .A(\myalu/myadder/myadder/c25 ), .Y(n923) );
  INVX1 U273 ( .A(\myalu/myadder/myadder/c21 ), .Y(n911) );
  INVX1 U274 ( .A(\myalu/myadder/myadder/c14 ), .Y(n890) );
  INVX1 U275 ( .A(\myalu/myadder/myadder/c18 ), .Y(n902) );
  INVX1 U276 ( .A(\myalu/myadder/myadder/c27 ), .Y(n929) );
  INVX1 U277 ( .A(\myalu/myadder/myadder/c28 ), .Y(n932) );
  INVX1 U278 ( .A(\myalu/myadder/myadder/c30 ), .Y(n938) );
  INVX1 U279 ( .A(\myalu/myadder/myadder/c29 ), .Y(n935) );
  INVX1 U280 ( .A(\myalu/myadder/myadder/c8 ), .Y(n872) );
  OR2X1 U281 ( .A(addr_b[2]), .B(n840), .Y(n194) );
  INVX1 U282 ( .A(n1042), .Y(\myalu/s0[9] ) );
  BUFX2 U283 ( .A(b[0]), .Y(n129) );
  INVX1 U284 ( .A(n311), .Y(n309) );
  INVX1 U285 ( .A(n311), .Y(n308) );
  INVX1 U286 ( .A(n311), .Y(n310) );
  INVX1 U287 ( .A(imm_en), .Y(n315) );
  INVX1 U288 ( .A(\myram/sel_s[0] ), .Y(n307) );
  INVX1 U289 ( .A(\myram/sel_s[8] ), .Y(n299) );
  INVX1 U290 ( .A(\myram/sel_s[2] ), .Y(n305) );
  INVX1 U291 ( .A(\myram/sel_s[6] ), .Y(n301) );
  INVX1 U292 ( .A(\myram/sel_s[7] ), .Y(n300) );
  INVX1 U293 ( .A(\myram/sel_s[10] ), .Y(n297) );
  INVX1 U294 ( .A(\myram/sel_s[11] ), .Y(n296) );
  INVX1 U295 ( .A(\myram/sel_s[15] ), .Y(n292) );
  INVX1 U296 ( .A(\myram/sel_s[1] ), .Y(n306) );
  INVX1 U297 ( .A(\myram/sel_s[5] ), .Y(n302) );
  INVX1 U298 ( .A(\myram/sel_s[9] ), .Y(n298) );
  INVX1 U299 ( .A(\myram/sel_s[13] ), .Y(n294) );
  AND2X1 U300 ( .A(alu_s[29]), .B(n315), .Y(mem_s[29]) );
  AND2X1 U301 ( .A(alu_s[26]), .B(n315), .Y(mem_s[26]) );
  AND2X1 U302 ( .A(alu_s[28]), .B(n315), .Y(mem_s[28]) );
  AND2X1 U303 ( .A(alu_s[18]), .B(n315), .Y(mem_s[18]) );
  AND2X1 U304 ( .A(alu_s[19]), .B(n315), .Y(mem_s[19]) );
  AND2X1 U305 ( .A(alu_s[20]), .B(n315), .Y(mem_s[20]) );
  AND2X1 U306 ( .A(alu_s[21]), .B(n315), .Y(mem_s[21]) );
  AND2X1 U307 ( .A(alu_s[22]), .B(n315), .Y(mem_s[22]) );
  AND2X1 U308 ( .A(alu_s[23]), .B(n315), .Y(mem_s[23]) );
  AND2X1 U309 ( .A(alu_s[24]), .B(n315), .Y(mem_s[24]) );
  AND2X1 U310 ( .A(alu_s[25]), .B(n315), .Y(mem_s[25]) );
  AND2X1 U311 ( .A(alu_s[27]), .B(n315), .Y(mem_s[27]) );
  INVX1 U312 ( .A(n235), .Y(n234) );
  INVX1 U313 ( .A(n219), .Y(n218) );
  INVX1 U314 ( .A(n291), .Y(n289) );
  INVX1 U315 ( .A(n227), .Y(n226) );
  INVX1 U316 ( .A(n243), .Y(n242) );
  INVX1 U317 ( .A(n239), .Y(n238) );
  INVX1 U318 ( .A(n237), .Y(n236) );
  INVX1 U319 ( .A(n231), .Y(n230) );
  INVX1 U320 ( .A(n229), .Y(n228) );
  INVX1 U321 ( .A(n223), .Y(n222) );
  INVX1 U322 ( .A(n221), .Y(n220) );
  INVX1 U323 ( .A(n215), .Y(n214) );
  INVX1 U324 ( .A(n213), .Y(n212) );
  INVX1 U325 ( .A(n241), .Y(n240) );
  INVX1 U326 ( .A(n233), .Y(n232) );
  INVX1 U327 ( .A(n225), .Y(n224) );
  INVX1 U328 ( .A(n217), .Y(n216) );
  INVX1 U329 ( .A(n1074), .Y(alu_s[9]) );
  AND2X1 U330 ( .A(alu_s[8]), .B(n315), .Y(mem_s[8]) );
  AND2X1 U331 ( .A(alu_s[10]), .B(n315), .Y(mem_s[10]) );
  AND2X1 U332 ( .A(alu_s[11]), .B(n315), .Y(mem_s[11]) );
  AND2X1 U333 ( .A(alu_s[12]), .B(n315), .Y(mem_s[12]) );
  AND2X1 U334 ( .A(alu_s[13]), .B(n315), .Y(mem_s[13]) );
  AND2X1 U335 ( .A(alu_s[14]), .B(n315), .Y(mem_s[14]) );
  AND2X1 U336 ( .A(alu_s[15]), .B(n315), .Y(mem_s[15]) );
  AND2X1 U337 ( .A(alu_s[16]), .B(n315), .Y(mem_s[16]) );
  AND2X1 U338 ( .A(alu_s[17]), .B(n315), .Y(mem_s[17]) );
  INVX1 U339 ( .A(n279), .Y(n278) );
  INVX1 U340 ( .A(n255), .Y(n254) );
  INVX1 U341 ( .A(n267), .Y(n266) );
  INVX1 U342 ( .A(n291), .Y(n290) );
  INVX1 U343 ( .A(n285), .Y(n284) );
  INVX1 U344 ( .A(n282), .Y(n281) );
  INVX1 U345 ( .A(n273), .Y(n272) );
  INVX1 U346 ( .A(n270), .Y(n269) );
  INVX1 U347 ( .A(n261), .Y(n260) );
  INVX1 U348 ( .A(n258), .Y(n257) );
  INVX1 U349 ( .A(n249), .Y(n248) );
  INVX1 U350 ( .A(n246), .Y(n245) );
  INVX1 U351 ( .A(n288), .Y(n287) );
  INVX1 U352 ( .A(n276), .Y(n275) );
  INVX1 U353 ( .A(n264), .Y(n263) );
  INVX1 U354 ( .A(n252), .Y(n251) );
  INVX1 U355 ( .A(alu_op[0]), .Y(n311) );
  INVX1 U356 ( .A(alu_op[2]), .Y(n314) );
  INVX1 U357 ( .A(n308), .Y(n312) );
  INVX1 U358 ( .A(\myram/sel_b[12] ), .Y(n255) );
  INVX1 U359 ( .A(\myram/sel_a[2] ), .Y(n239) );
  INVX1 U360 ( .A(\myram/sel_a[3] ), .Y(n237) );
  INVX1 U361 ( .A(\myram/sel_a[6] ), .Y(n231) );
  INVX1 U362 ( .A(\myram/sel_a[7] ), .Y(n229) );
  INVX1 U363 ( .A(\myram/sel_a[10] ), .Y(n223) );
  INVX1 U364 ( .A(\myram/sel_a[11] ), .Y(n221) );
  INVX1 U365 ( .A(\myram/sel_a[14] ), .Y(n215) );
  INVX1 U366 ( .A(\myram/sel_a[15] ), .Y(n213) );
  INVX1 U367 ( .A(\myram/sel_a[4] ), .Y(n235) );
  INVX1 U368 ( .A(\myram/sel_a[12] ), .Y(n219) );
  INVX1 U369 ( .A(\myram/sel_b[4] ), .Y(n279) );
  INVX1 U370 ( .A(\myram/sel_b[8] ), .Y(n267) );
  INVX1 U371 ( .A(\myram/sel_b[0] ), .Y(n291) );
  INVX1 U372 ( .A(\myram/sel_a[8] ), .Y(n227) );
  INVX1 U373 ( .A(\myram/sel_a[0] ), .Y(n243) );
  INVX1 U374 ( .A(\myram/sel_a[1] ), .Y(n241) );
  INVX1 U375 ( .A(\myram/sel_a[5] ), .Y(n233) );
  INVX1 U376 ( .A(\myram/sel_a[9] ), .Y(n225) );
  INVX1 U377 ( .A(\myram/sel_a[13] ), .Y(n217) );
  INVX1 U378 ( .A(\myram/sel_b[2] ), .Y(n285) );
  INVX1 U379 ( .A(\myram/sel_b[3] ), .Y(n282) );
  INVX1 U380 ( .A(\myram/sel_b[6] ), .Y(n273) );
  INVX1 U381 ( .A(\myram/sel_b[7] ), .Y(n270) );
  INVX1 U382 ( .A(\myram/sel_b[10] ), .Y(n261) );
  INVX1 U383 ( .A(\myram/sel_b[11] ), .Y(n258) );
  INVX1 U384 ( .A(\myram/sel_b[14] ), .Y(n249) );
  INVX1 U385 ( .A(\myram/sel_b[15] ), .Y(n246) );
  INVX1 U386 ( .A(\myram/sel_b[1] ), .Y(n288) );
  INVX1 U387 ( .A(\myram/sel_b[5] ), .Y(n276) );
  INVX1 U388 ( .A(\myram/sel_b[9] ), .Y(n264) );
  INVX1 U389 ( .A(\myram/sel_b[13] ), .Y(n252) );
  INVX1 U390 ( .A(n205), .Y(n833) );
  INVX1 U391 ( .A(n206), .Y(n832) );
  INVX1 U392 ( .A(n207), .Y(n829) );
  INVX1 U393 ( .A(n208), .Y(n828) );
  INVX1 U394 ( .A(n1062), .Y(\myalu/s0[29] ) );
  INVX1 U395 ( .A(n998), .Y(\myalu/s00[29] ) );
  INVX1 U396 ( .A(n1063), .Y(\myalu/s0[30] ) );
  INVX1 U397 ( .A(n999), .Y(\myalu/s00[30] ) );
  INVX1 U398 ( .A(n1064), .Y(\myalu/s0[31] ) );
  INVX1 U399 ( .A(n1000), .Y(\myalu/s00[31] ) );
  INVX1 U400 ( .A(n1051), .Y(\myalu/s0[18] ) );
  INVX1 U401 ( .A(n987), .Y(\myalu/s00[18] ) );
  INVX1 U402 ( .A(n1052), .Y(\myalu/s0[19] ) );
  INVX1 U403 ( .A(n988), .Y(\myalu/s00[19] ) );
  INVX1 U404 ( .A(n1053), .Y(\myalu/s0[20] ) );
  INVX1 U405 ( .A(n989), .Y(\myalu/s00[20] ) );
  INVX1 U406 ( .A(n1054), .Y(\myalu/s0[21] ) );
  INVX1 U407 ( .A(n990), .Y(\myalu/s00[21] ) );
  INVX1 U408 ( .A(n1055), .Y(\myalu/s0[22] ) );
  INVX1 U409 ( .A(n991), .Y(\myalu/s00[22] ) );
  INVX1 U410 ( .A(n1056), .Y(\myalu/s0[23] ) );
  INVX1 U411 ( .A(n992), .Y(\myalu/s00[23] ) );
  INVX1 U412 ( .A(n1057), .Y(\myalu/s0[24] ) );
  INVX1 U413 ( .A(n993), .Y(\myalu/s00[24] ) );
  INVX1 U414 ( .A(n1058), .Y(\myalu/s0[25] ) );
  INVX1 U415 ( .A(n994), .Y(\myalu/s00[25] ) );
  INVX1 U416 ( .A(n1059), .Y(\myalu/s0[26] ) );
  INVX1 U417 ( .A(n995), .Y(\myalu/s00[26] ) );
  INVX1 U418 ( .A(n1060), .Y(\myalu/s0[27] ) );
  INVX1 U419 ( .A(n996), .Y(\myalu/s00[27] ) );
  INVX1 U420 ( .A(n1061), .Y(\myalu/s0[28] ) );
  INVX1 U421 ( .A(n997), .Y(\myalu/s00[28] ) );
  INVX1 U422 ( .A(\alu_out/m0/n3 ), .Y(mem_s[0]) );
  INVX1 U423 ( .A(n1065), .Y(alu_s[0]) );
  INVX1 U424 ( .A(n943), .Y(mem_s[1]) );
  INVX1 U425 ( .A(n1066), .Y(alu_s[1]) );
  INVX1 U426 ( .A(n946), .Y(mem_s[4]) );
  INVX1 U427 ( .A(n1069), .Y(alu_s[4]) );
  INVX1 U428 ( .A(n947), .Y(mem_s[5]) );
  INVX1 U429 ( .A(n1070), .Y(alu_s[5]) );
  INVX1 U430 ( .A(n978), .Y(\myalu/s00[9] ) );
  AND2X1 U431 ( .A(\myalu/s10[9] ), .B(n313), .Y(n153) );
  INVX1 U432 ( .A(n1049), .Y(\myalu/s0[16] ) );
  INVX1 U433 ( .A(n985), .Y(\myalu/s00[16] ) );
  INVX1 U434 ( .A(n1050), .Y(\myalu/s0[17] ) );
  INVX1 U435 ( .A(n986), .Y(\myalu/s00[17] ) );
  INVX1 U436 ( .A(n1033), .Y(\myalu/s0[0] ) );
  INVX1 U437 ( .A(n969), .Y(\myalu/s00[0] ) );
  INVX1 U438 ( .A(n1034), .Y(\myalu/s0[1] ) );
  INVX1 U439 ( .A(n970), .Y(\myalu/s00[1] ) );
  INVX1 U440 ( .A(n1035), .Y(\myalu/s0[2] ) );
  INVX1 U441 ( .A(n971), .Y(\myalu/s00[2] ) );
  INVX1 U442 ( .A(n1036), .Y(\myalu/s0[3] ) );
  INVX1 U443 ( .A(n972), .Y(\myalu/s00[3] ) );
  INVX1 U444 ( .A(n1037), .Y(\myalu/s0[4] ) );
  INVX1 U445 ( .A(n973), .Y(\myalu/s00[4] ) );
  INVX1 U446 ( .A(n1038), .Y(\myalu/s0[5] ) );
  INVX1 U447 ( .A(n974), .Y(\myalu/s00[5] ) );
  INVX1 U448 ( .A(n1039), .Y(\myalu/s0[6] ) );
  INVX1 U449 ( .A(n975), .Y(\myalu/s00[6] ) );
  INVX1 U450 ( .A(n1040), .Y(\myalu/s0[7] ) );
  INVX1 U451 ( .A(n976), .Y(\myalu/s00[7] ) );
  INVX1 U452 ( .A(n1041), .Y(\myalu/s0[8] ) );
  INVX1 U453 ( .A(n977), .Y(\myalu/s00[8] ) );
  INVX1 U454 ( .A(n1043), .Y(\myalu/s0[10] ) );
  INVX1 U455 ( .A(n979), .Y(\myalu/s00[10] ) );
  INVX1 U456 ( .A(n1044), .Y(\myalu/s0[11] ) );
  INVX1 U457 ( .A(n980), .Y(\myalu/s00[11] ) );
  INVX1 U458 ( .A(n1045), .Y(\myalu/s0[12] ) );
  INVX1 U459 ( .A(n981), .Y(\myalu/s00[12] ) );
  INVX1 U460 ( .A(n1046), .Y(\myalu/s0[13] ) );
  INVX1 U461 ( .A(n982), .Y(\myalu/s00[13] ) );
  INVX1 U462 ( .A(n1047), .Y(\myalu/s0[14] ) );
  INVX1 U463 ( .A(n983), .Y(\myalu/s00[14] ) );
  INVX1 U464 ( .A(n1048), .Y(\myalu/s0[15] ) );
  INVX1 U465 ( .A(n984), .Y(\myalu/s00[15] ) );
  INVX1 U466 ( .A(n3), .Y(\mypc/branch_en ) );
  INVX1 U467 ( .A(n951), .Y(\mypc/temp_pc0[0] ) );
  INVX1 U468 ( .A(n953), .Y(\mypc/temp_pc0[1] ) );
  INVX1 U469 ( .A(\mypc/branch_en ), .Y(n952) );
  INVX1 U470 ( .A(n956), .Y(\mypc/temp_pc0[4] ) );
  INVX1 U471 ( .A(n957), .Y(\mypc/temp_pc0[5] ) );
  AND2X1 U472 ( .A(\myalu/s10[16] ), .B(n313), .Y(n154) );
  AND2X1 U473 ( .A(\myalu/s10[1] ), .B(n313), .Y(n155) );
  AND2X1 U474 ( .A(\myalu/s10[2] ), .B(n313), .Y(n156) );
  AND2X1 U475 ( .A(\myalu/s10[3] ), .B(n313), .Y(n157) );
  AND2X1 U476 ( .A(\myalu/s10[4] ), .B(n313), .Y(n158) );
  AND2X1 U477 ( .A(\myalu/s10[5] ), .B(n313), .Y(n159) );
  AND2X1 U478 ( .A(\myalu/s10[6] ), .B(n313), .Y(n160) );
  AND2X1 U479 ( .A(\myalu/s10[7] ), .B(n313), .Y(n161) );
  AND2X1 U480 ( .A(\myalu/s10[8] ), .B(n313), .Y(n162) );
  AND2X1 U481 ( .A(\myalu/s10[10] ), .B(n313), .Y(n163) );
  AND2X1 U482 ( .A(\myalu/s10[11] ), .B(n313), .Y(n164) );
  AND2X1 U483 ( .A(\myalu/s10[12] ), .B(n313), .Y(n165) );
  AND2X1 U484 ( .A(\myalu/s10[13] ), .B(n313), .Y(n166) );
  AND2X1 U485 ( .A(\myalu/s10[14] ), .B(n313), .Y(n167) );
  AND2X1 U486 ( .A(\myalu/s10[15] ), .B(n313), .Y(n168) );
  AND2X1 U487 ( .A(\myalu/s10[0] ), .B(n313), .Y(n169) );
  AND2X1 U488 ( .A(\myalu/s10[17] ), .B(n313), .Y(n170) );
  AND2X1 U489 ( .A(\myalu/s10[18] ), .B(n313), .Y(n171) );
  AND2X1 U490 ( .A(\myalu/s10[19] ), .B(n313), .Y(n172) );
  AND2X1 U491 ( .A(\myalu/s10[20] ), .B(n313), .Y(n173) );
  AND2X1 U492 ( .A(\myalu/s10[21] ), .B(n313), .Y(n174) );
  AND2X1 U493 ( .A(\myalu/s10[22] ), .B(n313), .Y(n175) );
  AND2X1 U494 ( .A(\myalu/s10[23] ), .B(n313), .Y(n176) );
  AND2X1 U495 ( .A(\myalu/s10[24] ), .B(n313), .Y(n177) );
  AND2X1 U496 ( .A(\myalu/s10[25] ), .B(n313), .Y(n178) );
  AND2X1 U497 ( .A(\myalu/s10[26] ), .B(n313), .Y(n179) );
  AND2X1 U498 ( .A(\myalu/s10[27] ), .B(n313), .Y(n180) );
  AND2X1 U499 ( .A(\myalu/s10[28] ), .B(n313), .Y(n181) );
  AND2X1 U500 ( .A(\myalu/s10[29] ), .B(n313), .Y(n182) );
  AND2X1 U501 ( .A(\myalu/s10[30] ), .B(n313), .Y(n183) );
  INVX1 U502 ( .A(n4), .Y(n2) );
  INVX1 U503 ( .A(\myram/sel_s[12] ), .Y(n295) );
  INVX1 U504 ( .A(\myram/sel_s[4] ), .Y(n303) );
  INVX1 U505 ( .A(\myram/sel_s[3] ), .Y(n304) );
  INVX1 U506 ( .A(\myram/sel_s[14] ), .Y(n293) );
  OR2X1 U507 ( .A(n843), .B(n186), .Y(n184) );
  INVX1 U508 ( .A(n209), .Y(n838) );
  INVX1 U509 ( .A(n211), .Y(n961) );
  INVX1 U510 ( .A(n210), .Y(n836) );
  AND2X1 U511 ( .A(\myalu/s10[31] ), .B(n313), .Y(n185) );
  OR2X1 U512 ( .A(n842), .B(\mypc/inc_pc[0] ), .Y(n186) );
  OR2X1 U513 ( .A(n844), .B(n184), .Y(n187) );
  OR2X1 U514 ( .A(n845), .B(n187), .Y(n188) );
  OR2X1 U515 ( .A(n846), .B(n188), .Y(n189) );
  OR2X1 U516 ( .A(n847), .B(n189), .Y(n190) );
  INVX1 U517 ( .A(alu_op[1]), .Y(n313) );
  BUFX2 U518 ( .A(addr_a[0]), .Y(n207) );
  BUFX2 U519 ( .A(addr_a[1]), .Y(n208) );
  OR2X1 U520 ( .A(addr_a[2]), .B(\myram/da/en0 ), .Y(n191) );
  OR2X1 U521 ( .A(addr_a[2]), .B(\myram/da/en1 ), .Y(n192) );
  OR2X1 U522 ( .A(addr_b[2]), .B(\myram/db/en1 ), .Y(n193) );
  INVX1 U523 ( .A(\myalu/myadder/myadder/c1 ), .Y(n851) );
  INVX1 U524 ( .A(\myram/db/d0/en1 ), .Y(n834) );
  AND2X1 U525 ( .A(addr_b[2]), .B(n840), .Y(\myram/db/d0/en1 ) );
  INVX1 U526 ( .A(\myram/da/d0/en1 ), .Y(n830) );
  AND2X1 U527 ( .A(addr_a[2]), .B(\myram/da/en0 ), .Y(\myram/da/d0/en1 ) );
  INVX1 U528 ( .A(\myram/da/d1/en1 ), .Y(n831) );
  AND2X1 U529 ( .A(addr_a[2]), .B(\myram/da/en1 ), .Y(\myram/da/d1/en1 ) );
  INVX1 U530 ( .A(\myalu/myadder/myadder/c31 ), .Y(n941) );
  INVX1 U531 ( .A(n1720), .Y(\myram/m1/mux_out[31] ) );
  INVX1 U532 ( .A(n1719), .Y(\myram/m1/mux_out[30] ) );
  INVX1 U533 ( .A(n1718), .Y(\myram/m1/mux_out[29] ) );
  INVX1 U534 ( .A(n1752), .Y(\myram/m2/mux_out[31] ) );
  INVX1 U535 ( .A(n1751), .Y(\myram/m2/mux_out[30] ) );
  INVX1 U536 ( .A(n1750), .Y(\myram/m2/mux_out[29] ) );
  INVX1 U537 ( .A(n1784), .Y(\myram/m3/mux_out[31] ) );
  INVX1 U538 ( .A(n1783), .Y(\myram/m3/mux_out[30] ) );
  INVX1 U539 ( .A(n1782), .Y(\myram/m3/mux_out[29] ) );
  INVX1 U540 ( .A(n1816), .Y(\myram/m4/mux_out[31] ) );
  INVX1 U541 ( .A(n1815), .Y(\myram/m4/mux_out[30] ) );
  INVX1 U542 ( .A(n1814), .Y(\myram/m4/mux_out[29] ) );
  INVX1 U543 ( .A(n1848), .Y(\myram/m5/mux_out[31] ) );
  INVX1 U544 ( .A(n1847), .Y(\myram/m5/mux_out[30] ) );
  INVX1 U545 ( .A(n1846), .Y(\myram/m5/mux_out[29] ) );
  INVX1 U546 ( .A(n1880), .Y(\myram/m6/mux_out[31] ) );
  INVX1 U547 ( .A(n1879), .Y(\myram/m6/mux_out[30] ) );
  INVX1 U548 ( .A(n1878), .Y(\myram/m6/mux_out[29] ) );
  INVX1 U549 ( .A(n1912), .Y(\myram/m7/mux_out[31] ) );
  INVX1 U550 ( .A(n1911), .Y(\myram/m7/mux_out[30] ) );
  INVX1 U551 ( .A(n1910), .Y(\myram/m7/mux_out[29] ) );
  INVX1 U552 ( .A(n1944), .Y(\myram/m8/mux_out[31] ) );
  INVX1 U553 ( .A(n1943), .Y(\myram/m8/mux_out[30] ) );
  INVX1 U554 ( .A(n1942), .Y(\myram/m8/mux_out[29] ) );
  INVX1 U555 ( .A(n1976), .Y(\myram/m9/mux_out[31] ) );
  INVX1 U556 ( .A(n1975), .Y(\myram/m9/mux_out[30] ) );
  INVX1 U557 ( .A(n1974), .Y(\myram/m9/mux_out[29] ) );
  INVX1 U558 ( .A(n2008), .Y(\myram/m10/mux_out[31] ) );
  INVX1 U559 ( .A(n2007), .Y(\myram/m10/mux_out[30] ) );
  INVX1 U560 ( .A(n2006), .Y(\myram/m10/mux_out[29] ) );
  INVX1 U561 ( .A(n2040), .Y(\myram/m11/mux_out[31] ) );
  INVX1 U562 ( .A(n2039), .Y(\myram/m11/mux_out[30] ) );
  INVX1 U563 ( .A(n2038), .Y(\myram/m11/mux_out[29] ) );
  INVX1 U564 ( .A(n2072), .Y(\myram/m12/mux_out[31] ) );
  INVX1 U565 ( .A(n2071), .Y(\myram/m12/mux_out[30] ) );
  INVX1 U566 ( .A(n2070), .Y(\myram/m12/mux_out[29] ) );
  INVX1 U567 ( .A(n2104), .Y(\myram/m13/mux_out[31] ) );
  INVX1 U568 ( .A(n2103), .Y(\myram/m13/mux_out[30] ) );
  INVX1 U569 ( .A(n2102), .Y(\myram/m13/mux_out[29] ) );
  INVX1 U570 ( .A(n2136), .Y(\myram/m14/mux_out[31] ) );
  INVX1 U571 ( .A(n2135), .Y(\myram/m14/mux_out[30] ) );
  INVX1 U572 ( .A(n2134), .Y(\myram/m14/mux_out[29] ) );
  INVX1 U573 ( .A(n2168), .Y(\myram/m15/mux_out[31] ) );
  INVX1 U574 ( .A(n2167), .Y(\myram/m15/mux_out[30] ) );
  INVX1 U575 ( .A(n2166), .Y(\myram/m15/mux_out[29] ) );
  INVX1 U576 ( .A(n1686), .Y(\myram/m0/mux_out[29] ) );
  INVX1 U577 ( .A(n1687), .Y(\myram/m0/mux_out[30] ) );
  INVX1 U578 ( .A(n1688), .Y(\myram/m0/mux_out[31] ) );
  INVX1 U579 ( .A(n1717), .Y(\myram/m1/mux_out[28] ) );
  INVX1 U580 ( .A(n1716), .Y(\myram/m1/mux_out[27] ) );
  INVX1 U581 ( .A(n1715), .Y(\myram/m1/mux_out[26] ) );
  INVX1 U582 ( .A(n1714), .Y(\myram/m1/mux_out[25] ) );
  INVX1 U583 ( .A(n1713), .Y(\myram/m1/mux_out[24] ) );
  INVX1 U584 ( .A(n1712), .Y(\myram/m1/mux_out[23] ) );
  INVX1 U585 ( .A(n1711), .Y(\myram/m1/mux_out[22] ) );
  INVX1 U586 ( .A(n1710), .Y(\myram/m1/mux_out[21] ) );
  INVX1 U587 ( .A(n1709), .Y(\myram/m1/mux_out[20] ) );
  INVX1 U588 ( .A(n1708), .Y(\myram/m1/mux_out[19] ) );
  INVX1 U589 ( .A(n1707), .Y(\myram/m1/mux_out[18] ) );
  INVX1 U590 ( .A(n1749), .Y(\myram/m2/mux_out[28] ) );
  INVX1 U591 ( .A(n1748), .Y(\myram/m2/mux_out[27] ) );
  INVX1 U592 ( .A(n1747), .Y(\myram/m2/mux_out[26] ) );
  INVX1 U593 ( .A(n1746), .Y(\myram/m2/mux_out[25] ) );
  INVX1 U594 ( .A(n1745), .Y(\myram/m2/mux_out[24] ) );
  INVX1 U595 ( .A(n1744), .Y(\myram/m2/mux_out[23] ) );
  INVX1 U596 ( .A(n1743), .Y(\myram/m2/mux_out[22] ) );
  INVX1 U597 ( .A(n1742), .Y(\myram/m2/mux_out[21] ) );
  INVX1 U598 ( .A(n1741), .Y(\myram/m2/mux_out[20] ) );
  INVX1 U599 ( .A(n1740), .Y(\myram/m2/mux_out[19] ) );
  INVX1 U600 ( .A(n1739), .Y(\myram/m2/mux_out[18] ) );
  INVX1 U601 ( .A(n1781), .Y(\myram/m3/mux_out[28] ) );
  INVX1 U602 ( .A(n1780), .Y(\myram/m3/mux_out[27] ) );
  INVX1 U603 ( .A(n1779), .Y(\myram/m3/mux_out[26] ) );
  INVX1 U604 ( .A(n1778), .Y(\myram/m3/mux_out[25] ) );
  INVX1 U605 ( .A(n1777), .Y(\myram/m3/mux_out[24] ) );
  INVX1 U606 ( .A(n1776), .Y(\myram/m3/mux_out[23] ) );
  INVX1 U607 ( .A(n1775), .Y(\myram/m3/mux_out[22] ) );
  INVX1 U608 ( .A(n1774), .Y(\myram/m3/mux_out[21] ) );
  INVX1 U609 ( .A(n1773), .Y(\myram/m3/mux_out[20] ) );
  INVX1 U610 ( .A(n1772), .Y(\myram/m3/mux_out[19] ) );
  INVX1 U611 ( .A(n1771), .Y(\myram/m3/mux_out[18] ) );
  INVX1 U612 ( .A(n1813), .Y(\myram/m4/mux_out[28] ) );
  INVX1 U613 ( .A(n1812), .Y(\myram/m4/mux_out[27] ) );
  INVX1 U614 ( .A(n1811), .Y(\myram/m4/mux_out[26] ) );
  INVX1 U615 ( .A(n1810), .Y(\myram/m4/mux_out[25] ) );
  INVX1 U616 ( .A(n1809), .Y(\myram/m4/mux_out[24] ) );
  INVX1 U617 ( .A(n1808), .Y(\myram/m4/mux_out[23] ) );
  INVX1 U618 ( .A(n1807), .Y(\myram/m4/mux_out[22] ) );
  INVX1 U619 ( .A(n1806), .Y(\myram/m4/mux_out[21] ) );
  INVX1 U620 ( .A(n1805), .Y(\myram/m4/mux_out[20] ) );
  INVX1 U621 ( .A(n1804), .Y(\myram/m4/mux_out[19] ) );
  INVX1 U622 ( .A(n1803), .Y(\myram/m4/mux_out[18] ) );
  INVX1 U623 ( .A(n1845), .Y(\myram/m5/mux_out[28] ) );
  INVX1 U624 ( .A(n1844), .Y(\myram/m5/mux_out[27] ) );
  INVX1 U625 ( .A(n1843), .Y(\myram/m5/mux_out[26] ) );
  INVX1 U626 ( .A(n1842), .Y(\myram/m5/mux_out[25] ) );
  INVX1 U627 ( .A(n1841), .Y(\myram/m5/mux_out[24] ) );
  INVX1 U628 ( .A(n1840), .Y(\myram/m5/mux_out[23] ) );
  INVX1 U629 ( .A(n1839), .Y(\myram/m5/mux_out[22] ) );
  INVX1 U630 ( .A(n1838), .Y(\myram/m5/mux_out[21] ) );
  INVX1 U631 ( .A(n1837), .Y(\myram/m5/mux_out[20] ) );
  INVX1 U632 ( .A(n1836), .Y(\myram/m5/mux_out[19] ) );
  INVX1 U633 ( .A(n1835), .Y(\myram/m5/mux_out[18] ) );
  INVX1 U634 ( .A(n1877), .Y(\myram/m6/mux_out[28] ) );
  INVX1 U635 ( .A(n1876), .Y(\myram/m6/mux_out[27] ) );
  INVX1 U636 ( .A(n1875), .Y(\myram/m6/mux_out[26] ) );
  INVX1 U637 ( .A(n1874), .Y(\myram/m6/mux_out[25] ) );
  INVX1 U638 ( .A(n1873), .Y(\myram/m6/mux_out[24] ) );
  INVX1 U639 ( .A(n1872), .Y(\myram/m6/mux_out[23] ) );
  INVX1 U640 ( .A(n1871), .Y(\myram/m6/mux_out[22] ) );
  INVX1 U641 ( .A(n1870), .Y(\myram/m6/mux_out[21] ) );
  INVX1 U642 ( .A(n1869), .Y(\myram/m6/mux_out[20] ) );
  INVX1 U643 ( .A(n1868), .Y(\myram/m6/mux_out[19] ) );
  INVX1 U644 ( .A(n1867), .Y(\myram/m6/mux_out[18] ) );
  INVX1 U645 ( .A(n1909), .Y(\myram/m7/mux_out[28] ) );
  INVX1 U646 ( .A(n1908), .Y(\myram/m7/mux_out[27] ) );
  INVX1 U647 ( .A(n1907), .Y(\myram/m7/mux_out[26] ) );
  INVX1 U648 ( .A(n1906), .Y(\myram/m7/mux_out[25] ) );
  INVX1 U649 ( .A(n1905), .Y(\myram/m7/mux_out[24] ) );
  INVX1 U650 ( .A(n1904), .Y(\myram/m7/mux_out[23] ) );
  INVX1 U651 ( .A(n1903), .Y(\myram/m7/mux_out[22] ) );
  INVX1 U652 ( .A(n1902), .Y(\myram/m7/mux_out[21] ) );
  INVX1 U653 ( .A(n1901), .Y(\myram/m7/mux_out[20] ) );
  INVX1 U654 ( .A(n1900), .Y(\myram/m7/mux_out[19] ) );
  INVX1 U655 ( .A(n1899), .Y(\myram/m7/mux_out[18] ) );
  INVX1 U656 ( .A(n1941), .Y(\myram/m8/mux_out[28] ) );
  INVX1 U657 ( .A(n1940), .Y(\myram/m8/mux_out[27] ) );
  INVX1 U658 ( .A(n1939), .Y(\myram/m8/mux_out[26] ) );
  INVX1 U659 ( .A(n1938), .Y(\myram/m8/mux_out[25] ) );
  INVX1 U660 ( .A(n1937), .Y(\myram/m8/mux_out[24] ) );
  INVX1 U661 ( .A(n1936), .Y(\myram/m8/mux_out[23] ) );
  INVX1 U662 ( .A(n1935), .Y(\myram/m8/mux_out[22] ) );
  INVX1 U663 ( .A(n1934), .Y(\myram/m8/mux_out[21] ) );
  INVX1 U664 ( .A(n1933), .Y(\myram/m8/mux_out[20] ) );
  INVX1 U665 ( .A(n1932), .Y(\myram/m8/mux_out[19] ) );
  INVX1 U666 ( .A(n1931), .Y(\myram/m8/mux_out[18] ) );
  INVX1 U667 ( .A(n1973), .Y(\myram/m9/mux_out[28] ) );
  INVX1 U668 ( .A(n1972), .Y(\myram/m9/mux_out[27] ) );
  INVX1 U669 ( .A(n1971), .Y(\myram/m9/mux_out[26] ) );
  INVX1 U670 ( .A(n1970), .Y(\myram/m9/mux_out[25] ) );
  INVX1 U671 ( .A(n1969), .Y(\myram/m9/mux_out[24] ) );
  INVX1 U672 ( .A(n1968), .Y(\myram/m9/mux_out[23] ) );
  INVX1 U673 ( .A(n1967), .Y(\myram/m9/mux_out[22] ) );
  INVX1 U674 ( .A(n1966), .Y(\myram/m9/mux_out[21] ) );
  INVX1 U675 ( .A(n1965), .Y(\myram/m9/mux_out[20] ) );
  INVX1 U676 ( .A(n1964), .Y(\myram/m9/mux_out[19] ) );
  INVX1 U677 ( .A(n1963), .Y(\myram/m9/mux_out[18] ) );
  INVX1 U678 ( .A(n2005), .Y(\myram/m10/mux_out[28] ) );
  INVX1 U679 ( .A(n2004), .Y(\myram/m10/mux_out[27] ) );
  INVX1 U680 ( .A(n2003), .Y(\myram/m10/mux_out[26] ) );
  INVX1 U681 ( .A(n2002), .Y(\myram/m10/mux_out[25] ) );
  INVX1 U682 ( .A(n2001), .Y(\myram/m10/mux_out[24] ) );
  INVX1 U683 ( .A(n2000), .Y(\myram/m10/mux_out[23] ) );
  INVX1 U684 ( .A(n1999), .Y(\myram/m10/mux_out[22] ) );
  INVX1 U685 ( .A(n1998), .Y(\myram/m10/mux_out[21] ) );
  INVX1 U686 ( .A(n1997), .Y(\myram/m10/mux_out[20] ) );
  INVX1 U687 ( .A(n1996), .Y(\myram/m10/mux_out[19] ) );
  INVX1 U688 ( .A(n1995), .Y(\myram/m10/mux_out[18] ) );
  INVX1 U689 ( .A(n2037), .Y(\myram/m11/mux_out[28] ) );
  INVX1 U690 ( .A(n2036), .Y(\myram/m11/mux_out[27] ) );
  INVX1 U691 ( .A(n2035), .Y(\myram/m11/mux_out[26] ) );
  INVX1 U692 ( .A(n2034), .Y(\myram/m11/mux_out[25] ) );
  INVX1 U693 ( .A(n2033), .Y(\myram/m11/mux_out[24] ) );
  INVX1 U694 ( .A(n2032), .Y(\myram/m11/mux_out[23] ) );
  INVX1 U695 ( .A(n2031), .Y(\myram/m11/mux_out[22] ) );
  INVX1 U696 ( .A(n2030), .Y(\myram/m11/mux_out[21] ) );
  INVX1 U697 ( .A(n2029), .Y(\myram/m11/mux_out[20] ) );
  INVX1 U698 ( .A(n2028), .Y(\myram/m11/mux_out[19] ) );
  INVX1 U699 ( .A(n2027), .Y(\myram/m11/mux_out[18] ) );
  INVX1 U700 ( .A(n2069), .Y(\myram/m12/mux_out[28] ) );
  INVX1 U701 ( .A(n2068), .Y(\myram/m12/mux_out[27] ) );
  INVX1 U702 ( .A(n2067), .Y(\myram/m12/mux_out[26] ) );
  INVX1 U703 ( .A(n2066), .Y(\myram/m12/mux_out[25] ) );
  INVX1 U704 ( .A(n2065), .Y(\myram/m12/mux_out[24] ) );
  INVX1 U705 ( .A(n2064), .Y(\myram/m12/mux_out[23] ) );
  INVX1 U706 ( .A(n2063), .Y(\myram/m12/mux_out[22] ) );
  INVX1 U707 ( .A(n2062), .Y(\myram/m12/mux_out[21] ) );
  INVX1 U708 ( .A(n2061), .Y(\myram/m12/mux_out[20] ) );
  INVX1 U709 ( .A(n2060), .Y(\myram/m12/mux_out[19] ) );
  INVX1 U710 ( .A(n2059), .Y(\myram/m12/mux_out[18] ) );
  INVX1 U711 ( .A(n2101), .Y(\myram/m13/mux_out[28] ) );
  INVX1 U712 ( .A(n2100), .Y(\myram/m13/mux_out[27] ) );
  INVX1 U713 ( .A(n2099), .Y(\myram/m13/mux_out[26] ) );
  INVX1 U714 ( .A(n2098), .Y(\myram/m13/mux_out[25] ) );
  INVX1 U715 ( .A(n2097), .Y(\myram/m13/mux_out[24] ) );
  INVX1 U716 ( .A(n2096), .Y(\myram/m13/mux_out[23] ) );
  INVX1 U717 ( .A(n2095), .Y(\myram/m13/mux_out[22] ) );
  INVX1 U718 ( .A(n2094), .Y(\myram/m13/mux_out[21] ) );
  INVX1 U719 ( .A(n2093), .Y(\myram/m13/mux_out[20] ) );
  INVX1 U720 ( .A(n2092), .Y(\myram/m13/mux_out[19] ) );
  INVX1 U721 ( .A(n2091), .Y(\myram/m13/mux_out[18] ) );
  INVX1 U722 ( .A(n2133), .Y(\myram/m14/mux_out[28] ) );
  INVX1 U723 ( .A(n2132), .Y(\myram/m14/mux_out[27] ) );
  INVX1 U724 ( .A(n2131), .Y(\myram/m14/mux_out[26] ) );
  INVX1 U725 ( .A(n2130), .Y(\myram/m14/mux_out[25] ) );
  INVX1 U726 ( .A(n2129), .Y(\myram/m14/mux_out[24] ) );
  INVX1 U727 ( .A(n2128), .Y(\myram/m14/mux_out[23] ) );
  INVX1 U728 ( .A(n2127), .Y(\myram/m14/mux_out[22] ) );
  INVX1 U729 ( .A(n2126), .Y(\myram/m14/mux_out[21] ) );
  INVX1 U730 ( .A(n2125), .Y(\myram/m14/mux_out[20] ) );
  INVX1 U731 ( .A(n2124), .Y(\myram/m14/mux_out[19] ) );
  INVX1 U732 ( .A(n2123), .Y(\myram/m14/mux_out[18] ) );
  INVX1 U733 ( .A(n2165), .Y(\myram/m15/mux_out[28] ) );
  INVX1 U734 ( .A(n2164), .Y(\myram/m15/mux_out[27] ) );
  INVX1 U735 ( .A(n2163), .Y(\myram/m15/mux_out[26] ) );
  INVX1 U736 ( .A(n2162), .Y(\myram/m15/mux_out[25] ) );
  INVX1 U737 ( .A(n2161), .Y(\myram/m15/mux_out[24] ) );
  INVX1 U738 ( .A(n2160), .Y(\myram/m15/mux_out[23] ) );
  INVX1 U739 ( .A(n2159), .Y(\myram/m15/mux_out[22] ) );
  INVX1 U740 ( .A(n2158), .Y(\myram/m15/mux_out[21] ) );
  INVX1 U741 ( .A(n2157), .Y(\myram/m15/mux_out[20] ) );
  INVX1 U742 ( .A(n2156), .Y(\myram/m15/mux_out[19] ) );
  INVX1 U743 ( .A(n2155), .Y(\myram/m15/mux_out[18] ) );
  INVX1 U744 ( .A(n1675), .Y(\myram/m0/mux_out[18] ) );
  INVX1 U745 ( .A(n1676), .Y(\myram/m0/mux_out[19] ) );
  INVX1 U746 ( .A(n1677), .Y(\myram/m0/mux_out[20] ) );
  INVX1 U747 ( .A(n1678), .Y(\myram/m0/mux_out[21] ) );
  INVX1 U748 ( .A(n1679), .Y(\myram/m0/mux_out[22] ) );
  INVX1 U749 ( .A(n1680), .Y(\myram/m0/mux_out[23] ) );
  INVX1 U750 ( .A(n1681), .Y(\myram/m0/mux_out[24] ) );
  INVX1 U751 ( .A(n1682), .Y(\myram/m0/mux_out[25] ) );
  INVX1 U752 ( .A(n1683), .Y(\myram/m0/mux_out[26] ) );
  INVX1 U753 ( .A(n1684), .Y(\myram/m0/mux_out[27] ) );
  INVX1 U754 ( .A(n1685), .Y(\myram/m0/mux_out[28] ) );
  INVX1 U755 ( .A(\myram/da/en1 ), .Y(\myram/da/en0 ) );
  INVX1 U756 ( .A(\myram/db/d1/en1 ), .Y(n835) );
  AND2X1 U757 ( .A(addr_b[2]), .B(\myram/db/en1 ), .Y(\myram/db/d1/en1 ) );
  INVX1 U758 ( .A(b[0]), .Y(n1416) );
  INVX1 U759 ( .A(b[0]), .Y(n1418) );
  INVX1 U760 ( .A(b[0]), .Y(n1157) );
  INVX1 U761 ( .A(n1421), .Y(\myalu/mysrl/s1[2] ) );
  INVX1 U762 ( .A(b[0]), .Y(n1420) );
  INVX1 U763 ( .A(n1423), .Y(\myalu/mysrl/s1[3] ) );
  INVX1 U764 ( .A(b[0]), .Y(n1422) );
  INVX1 U765 ( .A(n1425), .Y(\myalu/mysrl/s1[4] ) );
  INVX1 U766 ( .A(b[0]), .Y(n1424) );
  INVX1 U767 ( .A(n1427), .Y(\myalu/mysrl/s1[5] ) );
  INVX1 U768 ( .A(b[0]), .Y(n1426) );
  INVX1 U769 ( .A(n1429), .Y(\myalu/mysrl/s1[6] ) );
  INVX1 U770 ( .A(b[0]), .Y(n1428) );
  INVX1 U771 ( .A(n1430), .Y(\myalu/mysrl/s1[7] ) );
  INVX1 U772 ( .A(n1431), .Y(\myalu/mysrl/s1[8] ) );
  INVX1 U773 ( .A(n1432), .Y(\myalu/mysrl/s1[9] ) );
  INVX1 U774 ( .A(n1434), .Y(\myalu/mysrl/s1[10] ) );
  INVX1 U775 ( .A(b[0]), .Y(n1433) );
  INVX1 U776 ( .A(n1436), .Y(\myalu/mysrl/s1[11] ) );
  INVX1 U777 ( .A(b[0]), .Y(n1435) );
  INVX1 U778 ( .A(n1437), .Y(\myalu/mysrl/s1[12] ) );
  INVX1 U779 ( .A(n1438), .Y(\myalu/mysrl/s1[13] ) );
  INVX1 U780 ( .A(n1439), .Y(\myalu/mysrl/s1[14] ) );
  INVX1 U781 ( .A(n1441), .Y(\myalu/mysrl/s1[15] ) );
  INVX1 U782 ( .A(b[0]), .Y(n1440) );
  INVX1 U783 ( .A(n1442), .Y(\myalu/mysrl/s1[16] ) );
  INVX1 U784 ( .A(n1444), .Y(\myalu/mysrl/s1[17] ) );
  INVX1 U785 ( .A(b[0]), .Y(n1443) );
  INVX1 U786 ( .A(n1446), .Y(\myalu/mysrl/s1[18] ) );
  INVX1 U787 ( .A(b[0]), .Y(n1445) );
  INVX1 U788 ( .A(n1447), .Y(\myalu/mysrl/s1[19] ) );
  INVX1 U789 ( .A(n1448), .Y(\myalu/mysrl/s1[20] ) );
  INVX1 U790 ( .A(n1449), .Y(\myalu/mysrl/s1[21] ) );
  INVX1 U791 ( .A(n1451), .Y(\myalu/mysrl/s1[22] ) );
  INVX1 U792 ( .A(b[0]), .Y(n1450) );
  INVX1 U793 ( .A(n1452), .Y(\myalu/mysrl/s1[23] ) );
  INVX1 U794 ( .A(n1454), .Y(\myalu/mysrl/s1[24] ) );
  INVX1 U795 ( .A(b[0]), .Y(n1453) );
  INVX1 U796 ( .A(n1456), .Y(\myalu/mysrl/s1[25] ) );
  INVX1 U797 ( .A(b[0]), .Y(n1455) );
  INVX1 U798 ( .A(n1457), .Y(\myalu/mysrl/s1[26] ) );
  INVX1 U799 ( .A(n1458), .Y(\myalu/mysrl/s1[27] ) );
  INVX1 U800 ( .A(n1459), .Y(\myalu/mysrl/s1[28] ) );
  INVX1 U801 ( .A(n1461), .Y(\myalu/mysrl/s1[29] ) );
  INVX1 U802 ( .A(b[0]), .Y(n1460) );
  INVX1 U803 ( .A(n1114), .Y(\myalu/mysll/s1[8] ) );
  INVX1 U804 ( .A(b[0]), .Y(n1113) );
  INVX1 U805 ( .A(n1118), .Y(\myalu/mysll/s1[10] ) );
  INVX1 U806 ( .A(b[0]), .Y(n1117) );
  INVX1 U807 ( .A(n1122), .Y(\myalu/mysll/s1[12] ) );
  INVX1 U808 ( .A(b[0]), .Y(n1121) );
  INVX1 U809 ( .A(n1126), .Y(\myalu/mysll/s1[14] ) );
  INVX1 U810 ( .A(b[0]), .Y(n1125) );
  INVX1 U811 ( .A(n1106), .Y(\myalu/mysll/s1[4] ) );
  INVX1 U812 ( .A(b[0]), .Y(n1105) );
  INVX1 U813 ( .A(n1110), .Y(\myalu/mysll/s1[6] ) );
  INVX1 U814 ( .A(b[0]), .Y(n1109) );
  INVX1 U815 ( .A(n1102), .Y(\myalu/mysll/s1[2] ) );
  INVX1 U816 ( .A(b[0]), .Y(n1101) );
  INVX1 U817 ( .A(n1130), .Y(\myalu/mysll/s1[16] ) );
  INVX1 U818 ( .A(b[0]), .Y(n1129) );
  INVX1 U819 ( .A(n1134), .Y(\myalu/mysll/s1[18] ) );
  INVX1 U820 ( .A(b[0]), .Y(n1133) );
  INVX1 U821 ( .A(n1138), .Y(\myalu/mysll/s1[20] ) );
  INVX1 U822 ( .A(b[0]), .Y(n1137) );
  INVX1 U823 ( .A(n1142), .Y(\myalu/mysll/s1[22] ) );
  INVX1 U824 ( .A(b[0]), .Y(n1141) );
  INVX1 U825 ( .A(n1146), .Y(\myalu/mysll/s1[24] ) );
  INVX1 U826 ( .A(b[0]), .Y(n1145) );
  INVX1 U827 ( .A(n1150), .Y(\myalu/mysll/s1[26] ) );
  INVX1 U828 ( .A(b[0]), .Y(n1149) );
  INVX1 U829 ( .A(n1154), .Y(\myalu/mysll/s1[28] ) );
  INVX1 U830 ( .A(b[0]), .Y(n1153) );
  INVX1 U831 ( .A(n1462), .Y(\myalu/mysrl/s1[30] ) );
  INVX1 U832 ( .A(n1116), .Y(\myalu/mysll/s1[9] ) );
  INVX1 U833 ( .A(b[0]), .Y(n1115) );
  INVX1 U834 ( .A(n1120), .Y(\myalu/mysll/s1[11] ) );
  INVX1 U835 ( .A(b[0]), .Y(n1119) );
  INVX1 U836 ( .A(n1124), .Y(\myalu/mysll/s1[13] ) );
  INVX1 U837 ( .A(b[0]), .Y(n1123) );
  INVX1 U838 ( .A(n1128), .Y(\myalu/mysll/s1[15] ) );
  INVX1 U839 ( .A(b[0]), .Y(n1127) );
  INVX1 U840 ( .A(n1108), .Y(\myalu/mysll/s1[5] ) );
  INVX1 U841 ( .A(b[0]), .Y(n1107) );
  INVX1 U842 ( .A(n1112), .Y(\myalu/mysll/s1[7] ) );
  INVX1 U843 ( .A(b[0]), .Y(n1111) );
  INVX1 U844 ( .A(n1104), .Y(\myalu/mysll/s1[3] ) );
  INVX1 U845 ( .A(b[0]), .Y(n1103) );
  INVX1 U846 ( .A(n1100), .Y(\myalu/mysll/s1[1] ) );
  INVX1 U847 ( .A(b[0]), .Y(n1099) );
  INVX1 U848 ( .A(n1132), .Y(\myalu/mysll/s1[17] ) );
  INVX1 U849 ( .A(b[0]), .Y(n1131) );
  INVX1 U850 ( .A(n1136), .Y(\myalu/mysll/s1[19] ) );
  INVX1 U851 ( .A(b[0]), .Y(n1135) );
  INVX1 U852 ( .A(n1140), .Y(\myalu/mysll/s1[21] ) );
  INVX1 U853 ( .A(b[0]), .Y(n1139) );
  INVX1 U854 ( .A(n1144), .Y(\myalu/mysll/s1[23] ) );
  INVX1 U855 ( .A(b[0]), .Y(n1143) );
  INVX1 U856 ( .A(n1148), .Y(\myalu/mysll/s1[25] ) );
  INVX1 U857 ( .A(b[0]), .Y(n1147) );
  INVX1 U858 ( .A(n1152), .Y(\myalu/mysll/s1[27] ) );
  INVX1 U859 ( .A(b[0]), .Y(n1151) );
  INVX1 U860 ( .A(n1156), .Y(\myalu/mysll/s1[29] ) );
  INVX1 U861 ( .A(b[0]), .Y(n1155) );
  INVX1 U862 ( .A(n62), .Y(n1465) );
  INVX1 U863 ( .A(n1417), .Y(\myalu/mysrl/s1[0] ) );
  INVX1 U864 ( .A(n62), .Y(n1467) );
  INVX1 U865 ( .A(n1419), .Y(\myalu/mysrl/s1[1] ) );
  INVX1 U866 ( .A(n62), .Y(n1469) );
  INVX1 U867 ( .A(n62), .Y(n1471) );
  INVX1 U868 ( .A(n62), .Y(n1216) );
  INVX1 U869 ( .A(n62), .Y(n1218) );
  INVX1 U870 ( .A(n62), .Y(n1220) );
  INVX1 U871 ( .A(n1158), .Y(\myalu/mysll/s1[30] ) );
  INVX1 U872 ( .A(n62), .Y(n1222) );
  INVX1 U873 ( .A(n1159), .Y(\myalu/mysll/s1[31] ) );
  INVX1 U874 ( .A(n1474), .Y(\myalu/mysrl/s2[4] ) );
  INVX1 U875 ( .A(n62), .Y(n1473) );
  INVX1 U876 ( .A(n1476), .Y(\myalu/mysrl/s2[5] ) );
  INVX1 U877 ( .A(n62), .Y(n1475) );
  INVX1 U878 ( .A(n1477), .Y(\myalu/mysrl/s2[6] ) );
  INVX1 U879 ( .A(n1478), .Y(\myalu/mysrl/s2[7] ) );
  INVX1 U880 ( .A(n1480), .Y(\myalu/mysrl/s2[8] ) );
  INVX1 U881 ( .A(n62), .Y(n1479) );
  INVX1 U882 ( .A(n1481), .Y(\myalu/mysrl/s2[9] ) );
  INVX1 U883 ( .A(n1483), .Y(\myalu/mysrl/s2[10] ) );
  INVX1 U884 ( .A(n62), .Y(n1482) );
  INVX1 U885 ( .A(n1485), .Y(\myalu/mysrl/s2[11] ) );
  INVX1 U886 ( .A(n62), .Y(n1484) );
  INVX1 U887 ( .A(n1486), .Y(\myalu/mysrl/s2[12] ) );
  INVX1 U888 ( .A(n1487), .Y(\myalu/mysrl/s2[13] ) );
  INVX1 U889 ( .A(n1488), .Y(\myalu/mysrl/s2[14] ) );
  INVX1 U890 ( .A(n1489), .Y(\myalu/mysrl/s2[15] ) );
  INVX1 U891 ( .A(n1491), .Y(\myalu/mysrl/s2[16] ) );
  INVX1 U892 ( .A(n62), .Y(n1490) );
  INVX1 U893 ( .A(n1492), .Y(\myalu/mysrl/s2[17] ) );
  INVX1 U894 ( .A(n1494), .Y(\myalu/mysrl/s2[18] ) );
  INVX1 U895 ( .A(n62), .Y(n1493) );
  INVX1 U896 ( .A(n1496), .Y(\myalu/mysrl/s2[19] ) );
  INVX1 U897 ( .A(n62), .Y(n1495) );
  INVX1 U898 ( .A(n1498), .Y(\myalu/mysrl/s2[20] ) );
  INVX1 U899 ( .A(n62), .Y(n1497) );
  INVX1 U900 ( .A(n1499), .Y(\myalu/mysrl/s2[21] ) );
  INVX1 U901 ( .A(n1500), .Y(\myalu/mysrl/s2[22] ) );
  INVX1 U902 ( .A(n1501), .Y(\myalu/mysrl/s2[23] ) );
  INVX1 U903 ( .A(n1503), .Y(\myalu/mysrl/s2[24] ) );
  INVX1 U904 ( .A(n62), .Y(n1502) );
  INVX1 U905 ( .A(n1505), .Y(\myalu/mysrl/s2[25] ) );
  INVX1 U906 ( .A(n62), .Y(n1504) );
  INVX1 U907 ( .A(n1506), .Y(\myalu/mysrl/s2[26] ) );
  INVX1 U908 ( .A(n1507), .Y(\myalu/mysrl/s2[27] ) );
  INVX1 U909 ( .A(n1177), .Y(\myalu/mysll/s2[8] ) );
  INVX1 U910 ( .A(n62), .Y(n1176) );
  INVX1 U911 ( .A(n1185), .Y(\myalu/mysll/s2[12] ) );
  INVX1 U912 ( .A(n62), .Y(n1184) );
  INVX1 U913 ( .A(n1169), .Y(\myalu/mysll/s2[4] ) );
  INVX1 U914 ( .A(n62), .Y(n1168) );
  INVX1 U915 ( .A(n1193), .Y(\myalu/mysll/s2[16] ) );
  INVX1 U916 ( .A(n62), .Y(n1192) );
  INVX1 U917 ( .A(n1201), .Y(\myalu/mysll/s2[20] ) );
  INVX1 U918 ( .A(n62), .Y(n1200) );
  INVX1 U919 ( .A(n1209), .Y(\myalu/mysll/s2[24] ) );
  INVX1 U920 ( .A(n62), .Y(n1208) );
  INVX1 U921 ( .A(n1508), .Y(\myalu/mysrl/s2[28] ) );
  INVX1 U922 ( .A(n1179), .Y(\myalu/mysll/s2[9] ) );
  INVX1 U923 ( .A(n62), .Y(n1178) );
  INVX1 U924 ( .A(n1187), .Y(\myalu/mysll/s2[13] ) );
  INVX1 U925 ( .A(n62), .Y(n1186) );
  INVX1 U926 ( .A(n1171), .Y(\myalu/mysll/s2[5] ) );
  INVX1 U927 ( .A(n62), .Y(n1170) );
  INVX1 U928 ( .A(n1195), .Y(\myalu/mysll/s2[17] ) );
  INVX1 U929 ( .A(n62), .Y(n1194) );
  INVX1 U930 ( .A(n1203), .Y(\myalu/mysll/s2[21] ) );
  INVX1 U931 ( .A(n62), .Y(n1202) );
  INVX1 U932 ( .A(n1211), .Y(\myalu/mysll/s2[25] ) );
  INVX1 U933 ( .A(n62), .Y(n1210) );
  INVX1 U934 ( .A(n1510), .Y(\myalu/mysrl/s2[29] ) );
  INVX1 U935 ( .A(n62), .Y(n1509) );
  INVX1 U936 ( .A(n1181), .Y(\myalu/mysll/s2[10] ) );
  INVX1 U937 ( .A(n62), .Y(n1180) );
  INVX1 U938 ( .A(n1189), .Y(\myalu/mysll/s2[14] ) );
  INVX1 U939 ( .A(n62), .Y(n1188) );
  INVX1 U940 ( .A(n1173), .Y(\myalu/mysll/s2[6] ) );
  INVX1 U941 ( .A(n62), .Y(n1172) );
  INVX1 U942 ( .A(n1165), .Y(\myalu/mysll/s2[2] ) );
  INVX1 U943 ( .A(n62), .Y(n1164) );
  INVX1 U944 ( .A(n1197), .Y(\myalu/mysll/s2[18] ) );
  INVX1 U945 ( .A(n62), .Y(n1196) );
  INVX1 U946 ( .A(n1205), .Y(\myalu/mysll/s2[22] ) );
  INVX1 U947 ( .A(n62), .Y(n1204) );
  INVX1 U948 ( .A(n1213), .Y(\myalu/mysll/s2[26] ) );
  INVX1 U949 ( .A(n62), .Y(n1212) );
  INVX1 U950 ( .A(n1183), .Y(\myalu/mysll/s2[11] ) );
  INVX1 U951 ( .A(n62), .Y(n1182) );
  INVX1 U952 ( .A(n1191), .Y(\myalu/mysll/s2[15] ) );
  INVX1 U953 ( .A(n62), .Y(n1190) );
  INVX1 U954 ( .A(n1175), .Y(\myalu/mysll/s2[7] ) );
  INVX1 U955 ( .A(n62), .Y(n1174) );
  INVX1 U956 ( .A(n1167), .Y(\myalu/mysll/s2[3] ) );
  INVX1 U957 ( .A(n62), .Y(n1166) );
  INVX1 U958 ( .A(n1199), .Y(\myalu/mysll/s2[19] ) );
  INVX1 U959 ( .A(n62), .Y(n1198) );
  INVX1 U960 ( .A(n1207), .Y(\myalu/mysll/s2[23] ) );
  INVX1 U961 ( .A(n62), .Y(n1206) );
  INVX1 U962 ( .A(n1215), .Y(\myalu/mysll/s2[27] ) );
  INVX1 U963 ( .A(n62), .Y(n1214) );
  INVX1 U964 ( .A(n1527), .Y(\myalu/mysrl/s3[8] ) );
  INVX1 U965 ( .A(n25), .Y(n1526) );
  INVX1 U966 ( .A(n1529), .Y(\myalu/mysrl/s3[9] ) );
  INVX1 U967 ( .A(n25), .Y(n1528) );
  INVX1 U968 ( .A(n1531), .Y(\myalu/mysrl/s3[10] ) );
  INVX1 U969 ( .A(n25), .Y(n1530) );
  INVX1 U970 ( .A(n1533), .Y(\myalu/mysrl/s3[11] ) );
  INVX1 U971 ( .A(n25), .Y(n1532) );
  INVX1 U972 ( .A(n1535), .Y(\myalu/mysrl/s3[12] ) );
  INVX1 U973 ( .A(n25), .Y(n1534) );
  INVX1 U974 ( .A(n1536), .Y(\myalu/mysrl/s3[13] ) );
  INVX1 U975 ( .A(n1537), .Y(\myalu/mysrl/s3[14] ) );
  INVX1 U976 ( .A(n1538), .Y(\myalu/mysrl/s3[15] ) );
  INVX1 U977 ( .A(n1539), .Y(\myalu/mysrl/s3[16] ) );
  INVX1 U978 ( .A(n1540), .Y(\myalu/mysrl/s3[17] ) );
  INVX1 U979 ( .A(n1542), .Y(\myalu/mysrl/s3[18] ) );
  INVX1 U980 ( .A(n25), .Y(n1541) );
  INVX1 U981 ( .A(n1544), .Y(\myalu/mysrl/s3[19] ) );
  INVX1 U982 ( .A(n25), .Y(n1543) );
  INVX1 U983 ( .A(n1546), .Y(\myalu/mysrl/s3[20] ) );
  INVX1 U984 ( .A(n25), .Y(n1545) );
  INVX1 U985 ( .A(n1547), .Y(\myalu/mysrl/s3[21] ) );
  INVX1 U986 ( .A(n1548), .Y(\myalu/mysrl/s3[22] ) );
  INVX1 U987 ( .A(n1549), .Y(\myalu/mysrl/s3[23] ) );
  INVX1 U988 ( .A(n1257), .Y(\myalu/mysll/s3[16] ) );
  INVX1 U989 ( .A(n25), .Y(n1256) );
  INVX1 U990 ( .A(n1241), .Y(\myalu/mysll/s3[8] ) );
  INVX1 U991 ( .A(n25), .Y(n1240) );
  INVX1 U992 ( .A(n1551), .Y(\myalu/mysrl/s3[24] ) );
  INVX1 U993 ( .A(n25), .Y(n1550) );
  INVX1 U994 ( .A(n1259), .Y(\myalu/mysll/s3[17] ) );
  INVX1 U995 ( .A(n25), .Y(n1258) );
  INVX1 U996 ( .A(n1243), .Y(\myalu/mysll/s3[9] ) );
  INVX1 U997 ( .A(n25), .Y(n1242) );
  INVX1 U998 ( .A(n1553), .Y(\myalu/mysrl/s3[25] ) );
  INVX1 U999 ( .A(n25), .Y(n1552) );
  INVX1 U1000 ( .A(n1261), .Y(\myalu/mysll/s3[18] ) );
  INVX1 U1001 ( .A(n25), .Y(n1260) );
  INVX1 U1002 ( .A(n1245), .Y(\myalu/mysll/s3[10] ) );
  INVX1 U1003 ( .A(n25), .Y(n1244) );
  INVX1 U1004 ( .A(n1554), .Y(\myalu/mysrl/s3[26] ) );
  INVX1 U1005 ( .A(n1263), .Y(\myalu/mysll/s3[19] ) );
  INVX1 U1006 ( .A(n25), .Y(n1262) );
  INVX1 U1007 ( .A(n1247), .Y(\myalu/mysll/s3[11] ) );
  INVX1 U1008 ( .A(n25), .Y(n1246) );
  INVX1 U1009 ( .A(n1555), .Y(\myalu/mysrl/s3[27] ) );
  INVX1 U1010 ( .A(n1249), .Y(\myalu/mysll/s3[12] ) );
  INVX1 U1011 ( .A(n25), .Y(n1248) );
  INVX1 U1012 ( .A(n1233), .Y(\myalu/mysll/s3[4] ) );
  INVX1 U1013 ( .A(n25), .Y(n1232) );
  INVX1 U1014 ( .A(n1265), .Y(\myalu/mysll/s3[20] ) );
  INVX1 U1015 ( .A(n25), .Y(n1264) );
  INVX1 U1016 ( .A(n1251), .Y(\myalu/mysll/s3[13] ) );
  INVX1 U1017 ( .A(n25), .Y(n1250) );
  INVX1 U1018 ( .A(n1235), .Y(\myalu/mysll/s3[5] ) );
  INVX1 U1019 ( .A(n25), .Y(n1234) );
  INVX1 U1020 ( .A(n1267), .Y(\myalu/mysll/s3[21] ) );
  INVX1 U1021 ( .A(n25), .Y(n1266) );
  INVX1 U1022 ( .A(n1253), .Y(\myalu/mysll/s3[14] ) );
  INVX1 U1023 ( .A(n25), .Y(n1252) );
  INVX1 U1024 ( .A(n1237), .Y(\myalu/mysll/s3[6] ) );
  INVX1 U1025 ( .A(n25), .Y(n1236) );
  INVX1 U1026 ( .A(n1269), .Y(\myalu/mysll/s3[22] ) );
  INVX1 U1027 ( .A(n25), .Y(n1268) );
  INVX1 U1028 ( .A(n1255), .Y(\myalu/mysll/s3[15] ) );
  INVX1 U1029 ( .A(n25), .Y(n1254) );
  INVX1 U1030 ( .A(n1239), .Y(\myalu/mysll/s3[7] ) );
  INVX1 U1031 ( .A(n25), .Y(n1238) );
  INVX1 U1032 ( .A(n1271), .Y(\myalu/mysll/s3[23] ) );
  INVX1 U1033 ( .A(n25), .Y(n1270) );
  INVX1 U1034 ( .A(b[3]), .Y(n1576) );
  INVX1 U1035 ( .A(n1587), .Y(\myalu/mysrl/s4[16] ) );
  INVX1 U1036 ( .A(n1588), .Y(\myalu/mysrl/s4[17] ) );
  INVX1 U1037 ( .A(n1590), .Y(\myalu/mysrl/s4[18] ) );
  INVX1 U1038 ( .A(b[3]), .Y(n1589) );
  INVX1 U1039 ( .A(n1592), .Y(\myalu/mysrl/s4[19] ) );
  INVX1 U1040 ( .A(b[3]), .Y(n1591) );
  INVX1 U1041 ( .A(n1594), .Y(\myalu/mysrl/s4[20] ) );
  INVX1 U1042 ( .A(b[3]), .Y(n1593) );
  INVX1 U1043 ( .A(n1595), .Y(\myalu/mysrl/s4[21] ) );
  INVX1 U1044 ( .A(n1596), .Y(\myalu/mysrl/s4[22] ) );
  INVX1 U1045 ( .A(n1597), .Y(\myalu/mysrl/s4[23] ) );
  INVX1 U1046 ( .A(n1305), .Y(\myalu/mysll/s4[8] ) );
  INVX1 U1047 ( .A(b[3]), .Y(n1304) );
  INVX1 U1048 ( .A(n1307), .Y(\myalu/mysll/s4[9] ) );
  INVX1 U1049 ( .A(b[3]), .Y(n1306) );
  INVX1 U1050 ( .A(n1309), .Y(\myalu/mysll/s4[10] ) );
  INVX1 U1051 ( .A(b[3]), .Y(n1308) );
  INVX1 U1052 ( .A(n1311), .Y(\myalu/mysll/s4[11] ) );
  INVX1 U1053 ( .A(b[3]), .Y(n1310) );
  INVX1 U1054 ( .A(n1313), .Y(\myalu/mysll/s4[12] ) );
  INVX1 U1055 ( .A(b[3]), .Y(n1312) );
  INVX1 U1056 ( .A(n1315), .Y(\myalu/mysll/s4[13] ) );
  INVX1 U1057 ( .A(b[3]), .Y(n1314) );
  INVX1 U1058 ( .A(n1317), .Y(\myalu/mysll/s4[14] ) );
  INVX1 U1059 ( .A(b[3]), .Y(n1316) );
  INVX1 U1060 ( .A(n1319), .Y(\myalu/mysll/s4[15] ) );
  INVX1 U1061 ( .A(b[3]), .Y(n1318) );
  INVX1 U1062 ( .A(b[4]), .Y(n1609) );
  INVX1 U1063 ( .A(n1562), .Y(\myalu/mysrl/s4[0] ) );
  INVX1 U1064 ( .A(b[4]), .Y(n1611) );
  INVX1 U1065 ( .A(n1564), .Y(\myalu/mysrl/s4[1] ) );
  INVX1 U1066 ( .A(b[4]), .Y(n1613) );
  INVX1 U1067 ( .A(n1566), .Y(\myalu/mysrl/s4[2] ) );
  INVX1 U1068 ( .A(b[4]), .Y(n1615) );
  INVX1 U1069 ( .A(n1568), .Y(\myalu/mysrl/s4[3] ) );
  INVX1 U1070 ( .A(b[4]), .Y(n1617) );
  INVX1 U1071 ( .A(n1570), .Y(\myalu/mysrl/s4[4] ) );
  INVX1 U1072 ( .A(n1571), .Y(\myalu/mysrl/s4[5] ) );
  INVX1 U1073 ( .A(n1572), .Y(\myalu/mysrl/s4[6] ) );
  INVX1 U1074 ( .A(n1573), .Y(\myalu/mysrl/s4[7] ) );
  INVX1 U1075 ( .A(b[4]), .Y(n1622) );
  INVX1 U1076 ( .A(n1575), .Y(\myalu/mysrl/s4[8] ) );
  INVX1 U1077 ( .A(b[4]), .Y(n1626) );
  INVX1 U1078 ( .A(n1579), .Y(\myalu/mysrl/s4[10] ) );
  INVX1 U1079 ( .A(b[4]), .Y(n1628) );
  INVX1 U1080 ( .A(n1581), .Y(\myalu/mysrl/s4[11] ) );
  INVX1 U1081 ( .A(n1583), .Y(\myalu/mysrl/s4[12] ) );
  INVX1 U1082 ( .A(n1584), .Y(\myalu/mysrl/s4[13] ) );
  INVX1 U1083 ( .A(n1585), .Y(\myalu/mysrl/s4[14] ) );
  INVX1 U1084 ( .A(n1586), .Y(\myalu/mysrl/s4[15] ) );
  INVX1 U1085 ( .A(b[4]), .Y(n1384) );
  INVX1 U1086 ( .A(n1321), .Y(\myalu/mysll/s4[16] ) );
  INVX1 U1087 ( .A(b[4]), .Y(n1386) );
  INVX1 U1088 ( .A(n1323), .Y(\myalu/mysll/s4[17] ) );
  INVX1 U1089 ( .A(b[4]), .Y(n1388) );
  INVX1 U1090 ( .A(n1325), .Y(\myalu/mysll/s4[18] ) );
  INVX1 U1091 ( .A(b[4]), .Y(n1390) );
  INVX1 U1092 ( .A(n1327), .Y(\myalu/mysll/s4[19] ) );
  INVX1 U1093 ( .A(b[4]), .Y(n1392) );
  INVX1 U1094 ( .A(n1329), .Y(\myalu/mysll/s4[20] ) );
  INVX1 U1095 ( .A(b[4]), .Y(n1394) );
  INVX1 U1096 ( .A(n1331), .Y(\myalu/mysll/s4[21] ) );
  INVX1 U1097 ( .A(b[4]), .Y(n1396) );
  INVX1 U1098 ( .A(n1333), .Y(\myalu/mysll/s4[22] ) );
  INVX1 U1099 ( .A(b[4]), .Y(n1398) );
  INVX1 U1100 ( .A(n1335), .Y(\myalu/mysll/s4[23] ) );
  INVX1 U1101 ( .A(b[4]), .Y(n1400) );
  INVX1 U1102 ( .A(n1337), .Y(\myalu/mysll/s4[24] ) );
  INVX1 U1103 ( .A(b[4]), .Y(n1402) );
  INVX1 U1104 ( .A(n1339), .Y(\myalu/mysll/s4[25] ) );
  INVX1 U1105 ( .A(b[4]), .Y(n1404) );
  INVX1 U1106 ( .A(n1341), .Y(\myalu/mysll/s4[26] ) );
  INVX1 U1107 ( .A(b[4]), .Y(n1406) );
  INVX1 U1108 ( .A(n1343), .Y(\myalu/mysll/s4[27] ) );
  INVX1 U1109 ( .A(b[4]), .Y(n1408) );
  INVX1 U1110 ( .A(n1345), .Y(\myalu/mysll/s4[28] ) );
  INVX1 U1111 ( .A(b[4]), .Y(n1410) );
  INVX1 U1112 ( .A(n1347), .Y(\myalu/mysll/s4[29] ) );
  INVX1 U1113 ( .A(b[4]), .Y(n1412) );
  INVX1 U1114 ( .A(n1349), .Y(\myalu/mysll/s4[30] ) );
  INVX1 U1115 ( .A(b[4]), .Y(n1414) );
  INVX1 U1116 ( .A(n1351), .Y(\myalu/mysll/s4[31] ) );
  INVX1 U1117 ( .A(n1625), .Y(\myalu/ssr[9] ) );
  INVX1 U1118 ( .A(b[4]), .Y(n1624) );
  INVX1 U1119 ( .A(n1577), .Y(\myalu/mysrl/s4[9] ) );
  INVX1 U1120 ( .A(n1514), .Y(\myalu/mysrl/s3[0] ) );
  INVX1 U1121 ( .A(n25), .Y(n1513) );
  INVX1 U1122 ( .A(n1466), .Y(\myalu/mysrl/s2[0] ) );
  INVX1 U1123 ( .A(n1516), .Y(\myalu/mysrl/s3[1] ) );
  INVX1 U1124 ( .A(n25), .Y(n1515) );
  INVX1 U1125 ( .A(n1468), .Y(\myalu/mysrl/s2[1] ) );
  INVX1 U1126 ( .A(n1518), .Y(\myalu/mysrl/s3[2] ) );
  INVX1 U1127 ( .A(n25), .Y(n1517) );
  INVX1 U1128 ( .A(n1470), .Y(\myalu/mysrl/s2[2] ) );
  INVX1 U1129 ( .A(n1520), .Y(\myalu/mysrl/s3[3] ) );
  INVX1 U1130 ( .A(n25), .Y(n1519) );
  INVX1 U1131 ( .A(n1472), .Y(\myalu/mysrl/s2[3] ) );
  INVX1 U1132 ( .A(n1522), .Y(\myalu/mysrl/s3[4] ) );
  INVX1 U1133 ( .A(n25), .Y(n1521) );
  INVX1 U1134 ( .A(n1523), .Y(\myalu/mysrl/s3[5] ) );
  INVX1 U1135 ( .A(n1524), .Y(\myalu/mysrl/s3[6] ) );
  INVX1 U1136 ( .A(n1525), .Y(\myalu/mysrl/s3[7] ) );
  INVX1 U1137 ( .A(n1273), .Y(\myalu/mysll/s3[24] ) );
  INVX1 U1138 ( .A(n25), .Y(n1272) );
  INVX1 U1139 ( .A(n1275), .Y(\myalu/mysll/s3[25] ) );
  INVX1 U1140 ( .A(n25), .Y(n1274) );
  INVX1 U1141 ( .A(n1277), .Y(\myalu/mysll/s3[26] ) );
  INVX1 U1142 ( .A(n25), .Y(n1276) );
  INVX1 U1143 ( .A(n1279), .Y(\myalu/mysll/s3[27] ) );
  INVX1 U1144 ( .A(n25), .Y(n1278) );
  INVX1 U1145 ( .A(n1281), .Y(\myalu/mysll/s3[28] ) );
  INVX1 U1146 ( .A(n25), .Y(n1280) );
  INVX1 U1147 ( .A(n1217), .Y(\myalu/mysll/s2[28] ) );
  INVX1 U1148 ( .A(n1283), .Y(\myalu/mysll/s3[29] ) );
  INVX1 U1149 ( .A(n25), .Y(n1282) );
  INVX1 U1150 ( .A(n1219), .Y(\myalu/mysll/s2[29] ) );
  INVX1 U1151 ( .A(n1285), .Y(\myalu/mysll/s3[30] ) );
  INVX1 U1152 ( .A(n25), .Y(n1284) );
  INVX1 U1153 ( .A(n1221), .Y(\myalu/mysll/s2[30] ) );
  INVX1 U1154 ( .A(n1287), .Y(\myalu/mysll/s3[31] ) );
  INVX1 U1155 ( .A(n25), .Y(n1286) );
  INVX1 U1156 ( .A(n1223), .Y(\myalu/mysll/s2[31] ) );
  INVX1 U1157 ( .A(n944), .Y(mem_s[2]) );
  INVX1 U1158 ( .A(n1067), .Y(alu_s[2]) );
  INVX1 U1159 ( .A(n945), .Y(mem_s[3]) );
  INVX1 U1160 ( .A(n1068), .Y(alu_s[3]) );
  INVX1 U1161 ( .A(n948), .Y(mem_s[6]) );
  INVX1 U1162 ( .A(n1071), .Y(alu_s[6]) );
  INVX1 U1163 ( .A(n949), .Y(mem_s[7]) );
  INVX1 U1164 ( .A(n1072), .Y(alu_s[7]) );
  INVX1 U1165 ( .A(n1369), .Y(\myalu/ssl[8] ) );
  INVX1 U1166 ( .A(n1623), .Y(\myalu/ssr[8] ) );
  INVX1 U1167 ( .A(n1373), .Y(\myalu/ssl[10] ) );
  INVX1 U1168 ( .A(n1627), .Y(\myalu/ssr[10] ) );
  INVX1 U1169 ( .A(n1375), .Y(\myalu/ssl[11] ) );
  INVX1 U1170 ( .A(n1629), .Y(\myalu/ssr[11] ) );
  INVX1 U1171 ( .A(n1377), .Y(\myalu/ssl[12] ) );
  INVX1 U1172 ( .A(n1630), .Y(\myalu/ssr[12] ) );
  INVX1 U1173 ( .A(n1379), .Y(\myalu/ssl[13] ) );
  INVX1 U1174 ( .A(n1631), .Y(\myalu/ssr[13] ) );
  INVX1 U1175 ( .A(n1381), .Y(\myalu/ssl[14] ) );
  INVX1 U1176 ( .A(n1632), .Y(\myalu/ssr[14] ) );
  INVX1 U1177 ( .A(n1383), .Y(\myalu/ssl[15] ) );
  INVX1 U1178 ( .A(n1633), .Y(\myalu/ssr[15] ) );
  INVX1 U1179 ( .A(n1353), .Y(\myalu/ssl[0] ) );
  INVX1 U1180 ( .A(n1610), .Y(\myalu/ssr[0] ) );
  INVX1 U1181 ( .A(n1355), .Y(\myalu/ssl[1] ) );
  INVX1 U1182 ( .A(n1612), .Y(\myalu/ssr[1] ) );
  INVX1 U1183 ( .A(n1357), .Y(\myalu/ssl[2] ) );
  INVX1 U1184 ( .A(n1614), .Y(\myalu/ssr[2] ) );
  INVX1 U1185 ( .A(n1359), .Y(\myalu/ssl[3] ) );
  INVX1 U1186 ( .A(n1616), .Y(\myalu/ssr[3] ) );
  INVX1 U1187 ( .A(n1361), .Y(\myalu/ssl[4] ) );
  INVX1 U1188 ( .A(n1618), .Y(\myalu/ssr[4] ) );
  INVX1 U1189 ( .A(n1363), .Y(\myalu/ssl[5] ) );
  INVX1 U1190 ( .A(n1619), .Y(\myalu/ssr[5] ) );
  INVX1 U1191 ( .A(n1365), .Y(\myalu/ssl[6] ) );
  INVX1 U1192 ( .A(n1620), .Y(\myalu/ssr[6] ) );
  INVX1 U1193 ( .A(n1367), .Y(\myalu/ssl[7] ) );
  INVX1 U1194 ( .A(n1621), .Y(\myalu/ssr[7] ) );
  INVX1 U1195 ( .A(n1225), .Y(\myalu/mysll/s3[0] ) );
  INVX1 U1196 ( .A(n25), .Y(n1224) );
  INVX1 U1197 ( .A(n1635), .Y(\myalu/ssr[16] ) );
  INVX1 U1198 ( .A(n1385), .Y(\myalu/ssl[16] ) );
  INVX1 U1199 ( .A(n1637), .Y(\myalu/ssr[17] ) );
  INVX1 U1200 ( .A(n1387), .Y(\myalu/ssl[17] ) );
  INVX1 U1201 ( .A(n1639), .Y(\myalu/ssr[18] ) );
  INVX1 U1202 ( .A(n1389), .Y(\myalu/ssl[18] ) );
  INVX1 U1203 ( .A(n1641), .Y(\myalu/ssr[19] ) );
  INVX1 U1204 ( .A(n1391), .Y(\myalu/ssl[19] ) );
  INVX1 U1205 ( .A(n1643), .Y(\myalu/ssr[20] ) );
  INVX1 U1206 ( .A(n1393), .Y(\myalu/ssl[20] ) );
  INVX1 U1207 ( .A(n1644), .Y(\myalu/ssr[21] ) );
  INVX1 U1208 ( .A(n1395), .Y(\myalu/ssl[21] ) );
  INVX1 U1209 ( .A(n1645), .Y(\myalu/ssr[22] ) );
  INVX1 U1210 ( .A(n1397), .Y(\myalu/ssl[22] ) );
  INVX1 U1211 ( .A(n1646), .Y(\myalu/ssr[23] ) );
  INVX1 U1212 ( .A(n1399), .Y(\myalu/ssl[23] ) );
  INVX1 U1213 ( .A(n1648), .Y(\myalu/ssr[24] ) );
  INVX1 U1214 ( .A(n1401), .Y(\myalu/ssl[24] ) );
  INVX1 U1215 ( .A(n1649), .Y(\myalu/ssr[25] ) );
  INVX1 U1216 ( .A(n1403), .Y(\myalu/ssl[25] ) );
  INVX1 U1217 ( .A(n1651), .Y(\myalu/ssr[26] ) );
  INVX1 U1218 ( .A(n1405), .Y(\myalu/ssl[26] ) );
  INVX1 U1219 ( .A(n1652), .Y(\myalu/ssr[27] ) );
  INVX1 U1220 ( .A(n1407), .Y(\myalu/ssl[27] ) );
  INVX1 U1221 ( .A(n1653), .Y(\myalu/ssr[28] ) );
  INVX1 U1222 ( .A(n1409), .Y(\myalu/ssl[28] ) );
  INVX1 U1223 ( .A(n1654), .Y(\myalu/ssr[29] ) );
  INVX1 U1224 ( .A(n1411), .Y(\myalu/ssl[29] ) );
  INVX1 U1225 ( .A(n1655), .Y(\myalu/ssr[30] ) );
  INVX1 U1226 ( .A(n1413), .Y(\myalu/ssl[30] ) );
  INVX1 U1227 ( .A(n1656), .Y(\myalu/ssr[31] ) );
  INVX1 U1228 ( .A(n1415), .Y(\myalu/ssl[31] ) );
  INVX1 U1229 ( .A(n1161), .Y(\myalu/mysll/s2[0] ) );
  INVX1 U1230 ( .A(n62), .Y(n1160) );
  INVX1 U1231 ( .A(n1227), .Y(\myalu/mysll/s3[1] ) );
  INVX1 U1232 ( .A(n25), .Y(n1226) );
  INVX1 U1233 ( .A(n1559), .Y(\myalu/mysrl/s3[30] ) );
  INVX1 U1234 ( .A(n1293), .Y(\myalu/mysll/s4[2] ) );
  INVX1 U1235 ( .A(b[3]), .Y(n1292) );
  INVX1 U1236 ( .A(n1295), .Y(\myalu/mysll/s4[3] ) );
  INVX1 U1237 ( .A(b[3]), .Y(n1294) );
  INVX1 U1238 ( .A(n1605), .Y(\myalu/mysrl/s4[28] ) );
  INVX1 U1239 ( .A(b[3]), .Y(n1604) );
  INVX1 U1240 ( .A(n1606), .Y(\myalu/mysrl/s4[29] ) );
  INVX1 U1241 ( .A(n1289), .Y(\myalu/mysll/s4[0] ) );
  INVX1 U1242 ( .A(b[3]), .Y(n1288) );
  INVX1 U1243 ( .A(n1291), .Y(\myalu/mysll/s4[1] ) );
  INVX1 U1244 ( .A(b[3]), .Y(n1290) );
  INVX1 U1245 ( .A(n1607), .Y(\myalu/mysrl/s4[30] ) );
  INVX1 U1246 ( .A(n1098), .Y(\myalu/mysll/s1[0] ) );
  INVX1 U1247 ( .A(b[0]), .Y(n1097) );
  INVX1 U1248 ( .A(n1163), .Y(\myalu/mysll/s2[1] ) );
  INVX1 U1249 ( .A(n62), .Y(n1162) );
  INVX1 U1250 ( .A(n1511), .Y(\myalu/mysrl/s2[30] ) );
  INVX1 U1251 ( .A(n1229), .Y(\myalu/mysll/s3[2] ) );
  INVX1 U1252 ( .A(n25), .Y(n1228) );
  INVX1 U1253 ( .A(n1231), .Y(\myalu/mysll/s3[3] ) );
  INVX1 U1254 ( .A(n25), .Y(n1230) );
  INVX1 U1255 ( .A(n1557), .Y(\myalu/mysrl/s3[28] ) );
  INVX1 U1256 ( .A(n25), .Y(n1556) );
  INVX1 U1257 ( .A(n1558), .Y(\myalu/mysrl/s3[29] ) );
  INVX1 U1258 ( .A(n1297), .Y(\myalu/mysll/s4[4] ) );
  INVX1 U1259 ( .A(b[3]), .Y(n1296) );
  INVX1 U1260 ( .A(n1299), .Y(\myalu/mysll/s4[5] ) );
  INVX1 U1261 ( .A(b[3]), .Y(n1298) );
  INVX1 U1262 ( .A(n1301), .Y(\myalu/mysll/s4[6] ) );
  INVX1 U1263 ( .A(b[3]), .Y(n1300) );
  INVX1 U1264 ( .A(n1303), .Y(\myalu/mysll/s4[7] ) );
  INVX1 U1265 ( .A(b[3]), .Y(n1302) );
  INVX1 U1266 ( .A(n1599), .Y(\myalu/mysrl/s4[24] ) );
  INVX1 U1267 ( .A(b[3]), .Y(n1598) );
  INVX1 U1268 ( .A(n1601), .Y(\myalu/mysrl/s4[25] ) );
  INVX1 U1269 ( .A(b[3]), .Y(n1600) );
  INVX1 U1270 ( .A(n1602), .Y(\myalu/mysrl/s4[26] ) );
  INVX1 U1271 ( .A(n1603), .Y(\myalu/mysrl/s4[27] ) );
  INVX1 U1272 ( .A(n1371), .Y(\myalu/ssl[9] ) );
  INVX1 U1273 ( .A(b[4]), .Y(n1370) );
  INVX1 U1274 ( .A(n1706), .Y(\myram/m1/mux_out[17] ) );
  INVX1 U1275 ( .A(n1705), .Y(\myram/m1/mux_out[16] ) );
  INVX1 U1276 ( .A(n1704), .Y(\myram/m1/mux_out[15] ) );
  INVX1 U1277 ( .A(n1703), .Y(\myram/m1/mux_out[14] ) );
  INVX1 U1278 ( .A(n1702), .Y(\myram/m1/mux_out[13] ) );
  INVX1 U1279 ( .A(n1701), .Y(\myram/m1/mux_out[12] ) );
  INVX1 U1280 ( .A(n1700), .Y(\myram/m1/mux_out[11] ) );
  INVX1 U1281 ( .A(n1699), .Y(\myram/m1/mux_out[10] ) );
  INVX1 U1282 ( .A(n1698), .Y(\myram/m1/mux_out[9] ) );
  INVX1 U1283 ( .A(n1697), .Y(\myram/m1/mux_out[8] ) );
  INVX1 U1284 ( .A(n1696), .Y(\myram/m1/mux_out[7] ) );
  INVX1 U1285 ( .A(n1695), .Y(\myram/m1/mux_out[6] ) );
  INVX1 U1286 ( .A(n1694), .Y(\myram/m1/mux_out[5] ) );
  INVX1 U1287 ( .A(n1693), .Y(\myram/m1/mux_out[4] ) );
  INVX1 U1288 ( .A(n1692), .Y(\myram/m1/mux_out[3] ) );
  INVX1 U1289 ( .A(n1691), .Y(\myram/m1/mux_out[2] ) );
  INVX1 U1290 ( .A(n1690), .Y(\myram/m1/mux_out[1] ) );
  INVX1 U1291 ( .A(n1689), .Y(\myram/m1/mux_out[0] ) );
  INVX1 U1292 ( .A(n1738), .Y(\myram/m2/mux_out[17] ) );
  INVX1 U1293 ( .A(n1737), .Y(\myram/m2/mux_out[16] ) );
  INVX1 U1294 ( .A(n1736), .Y(\myram/m2/mux_out[15] ) );
  INVX1 U1295 ( .A(n1735), .Y(\myram/m2/mux_out[14] ) );
  INVX1 U1296 ( .A(n1734), .Y(\myram/m2/mux_out[13] ) );
  INVX1 U1297 ( .A(n1733), .Y(\myram/m2/mux_out[12] ) );
  INVX1 U1298 ( .A(n1732), .Y(\myram/m2/mux_out[11] ) );
  INVX1 U1299 ( .A(n1731), .Y(\myram/m2/mux_out[10] ) );
  INVX1 U1300 ( .A(n1730), .Y(\myram/m2/mux_out[9] ) );
  INVX1 U1301 ( .A(n1729), .Y(\myram/m2/mux_out[8] ) );
  INVX1 U1302 ( .A(n1728), .Y(\myram/m2/mux_out[7] ) );
  INVX1 U1303 ( .A(n1727), .Y(\myram/m2/mux_out[6] ) );
  INVX1 U1304 ( .A(n1726), .Y(\myram/m2/mux_out[5] ) );
  INVX1 U1305 ( .A(n1725), .Y(\myram/m2/mux_out[4] ) );
  INVX1 U1306 ( .A(n1724), .Y(\myram/m2/mux_out[3] ) );
  INVX1 U1307 ( .A(n1723), .Y(\myram/m2/mux_out[2] ) );
  INVX1 U1308 ( .A(n1722), .Y(\myram/m2/mux_out[1] ) );
  INVX1 U1309 ( .A(n1721), .Y(\myram/m2/mux_out[0] ) );
  INVX1 U1310 ( .A(n1770), .Y(\myram/m3/mux_out[17] ) );
  INVX1 U1311 ( .A(n1769), .Y(\myram/m3/mux_out[16] ) );
  INVX1 U1312 ( .A(n1768), .Y(\myram/m3/mux_out[15] ) );
  INVX1 U1313 ( .A(n1767), .Y(\myram/m3/mux_out[14] ) );
  INVX1 U1314 ( .A(n1766), .Y(\myram/m3/mux_out[13] ) );
  INVX1 U1315 ( .A(n1765), .Y(\myram/m3/mux_out[12] ) );
  INVX1 U1316 ( .A(n1764), .Y(\myram/m3/mux_out[11] ) );
  INVX1 U1317 ( .A(n1763), .Y(\myram/m3/mux_out[10] ) );
  INVX1 U1318 ( .A(n1762), .Y(\myram/m3/mux_out[9] ) );
  INVX1 U1319 ( .A(n1761), .Y(\myram/m3/mux_out[8] ) );
  INVX1 U1320 ( .A(n1760), .Y(\myram/m3/mux_out[7] ) );
  INVX1 U1321 ( .A(n1759), .Y(\myram/m3/mux_out[6] ) );
  INVX1 U1322 ( .A(n1758), .Y(\myram/m3/mux_out[5] ) );
  INVX1 U1323 ( .A(n1757), .Y(\myram/m3/mux_out[4] ) );
  INVX1 U1324 ( .A(n1756), .Y(\myram/m3/mux_out[3] ) );
  INVX1 U1325 ( .A(n1755), .Y(\myram/m3/mux_out[2] ) );
  INVX1 U1326 ( .A(n1754), .Y(\myram/m3/mux_out[1] ) );
  INVX1 U1327 ( .A(n1753), .Y(\myram/m3/mux_out[0] ) );
  INVX1 U1328 ( .A(n1802), .Y(\myram/m4/mux_out[17] ) );
  INVX1 U1329 ( .A(n1801), .Y(\myram/m4/mux_out[16] ) );
  INVX1 U1330 ( .A(n1800), .Y(\myram/m4/mux_out[15] ) );
  INVX1 U1331 ( .A(n1799), .Y(\myram/m4/mux_out[14] ) );
  INVX1 U1332 ( .A(n1798), .Y(\myram/m4/mux_out[13] ) );
  INVX1 U1333 ( .A(n1797), .Y(\myram/m4/mux_out[12] ) );
  INVX1 U1334 ( .A(n1796), .Y(\myram/m4/mux_out[11] ) );
  INVX1 U1335 ( .A(n1795), .Y(\myram/m4/mux_out[10] ) );
  INVX1 U1336 ( .A(n1794), .Y(\myram/m4/mux_out[9] ) );
  INVX1 U1337 ( .A(n1793), .Y(\myram/m4/mux_out[8] ) );
  INVX1 U1338 ( .A(n1792), .Y(\myram/m4/mux_out[7] ) );
  INVX1 U1339 ( .A(n1791), .Y(\myram/m4/mux_out[6] ) );
  INVX1 U1340 ( .A(n1790), .Y(\myram/m4/mux_out[5] ) );
  INVX1 U1341 ( .A(n1789), .Y(\myram/m4/mux_out[4] ) );
  INVX1 U1342 ( .A(n1788), .Y(\myram/m4/mux_out[3] ) );
  INVX1 U1343 ( .A(n1787), .Y(\myram/m4/mux_out[2] ) );
  INVX1 U1344 ( .A(n1786), .Y(\myram/m4/mux_out[1] ) );
  INVX1 U1345 ( .A(n1785), .Y(\myram/m4/mux_out[0] ) );
  INVX1 U1346 ( .A(n1834), .Y(\myram/m5/mux_out[17] ) );
  INVX1 U1347 ( .A(n1833), .Y(\myram/m5/mux_out[16] ) );
  INVX1 U1348 ( .A(n1832), .Y(\myram/m5/mux_out[15] ) );
  INVX1 U1349 ( .A(n1831), .Y(\myram/m5/mux_out[14] ) );
  INVX1 U1350 ( .A(n1830), .Y(\myram/m5/mux_out[13] ) );
  INVX1 U1351 ( .A(n1829), .Y(\myram/m5/mux_out[12] ) );
  INVX1 U1352 ( .A(n1828), .Y(\myram/m5/mux_out[11] ) );
  INVX1 U1353 ( .A(n1827), .Y(\myram/m5/mux_out[10] ) );
  INVX1 U1354 ( .A(n1826), .Y(\myram/m5/mux_out[9] ) );
  INVX1 U1355 ( .A(n1825), .Y(\myram/m5/mux_out[8] ) );
  INVX1 U1356 ( .A(n1824), .Y(\myram/m5/mux_out[7] ) );
  INVX1 U1357 ( .A(n1823), .Y(\myram/m5/mux_out[6] ) );
  INVX1 U1358 ( .A(n1822), .Y(\myram/m5/mux_out[5] ) );
  INVX1 U1359 ( .A(n1821), .Y(\myram/m5/mux_out[4] ) );
  INVX1 U1360 ( .A(n1820), .Y(\myram/m5/mux_out[3] ) );
  INVX1 U1361 ( .A(n1819), .Y(\myram/m5/mux_out[2] ) );
  INVX1 U1362 ( .A(n1818), .Y(\myram/m5/mux_out[1] ) );
  INVX1 U1363 ( .A(n1817), .Y(\myram/m5/mux_out[0] ) );
  INVX1 U1364 ( .A(n1866), .Y(\myram/m6/mux_out[17] ) );
  INVX1 U1365 ( .A(n1865), .Y(\myram/m6/mux_out[16] ) );
  INVX1 U1366 ( .A(n1864), .Y(\myram/m6/mux_out[15] ) );
  INVX1 U1367 ( .A(n1863), .Y(\myram/m6/mux_out[14] ) );
  INVX1 U1368 ( .A(n1862), .Y(\myram/m6/mux_out[13] ) );
  INVX1 U1369 ( .A(n1861), .Y(\myram/m6/mux_out[12] ) );
  INVX1 U1370 ( .A(n1860), .Y(\myram/m6/mux_out[11] ) );
  INVX1 U1371 ( .A(n1859), .Y(\myram/m6/mux_out[10] ) );
  INVX1 U1372 ( .A(n1858), .Y(\myram/m6/mux_out[9] ) );
  INVX1 U1373 ( .A(n1857), .Y(\myram/m6/mux_out[8] ) );
  INVX1 U1374 ( .A(n1856), .Y(\myram/m6/mux_out[7] ) );
  INVX1 U1375 ( .A(n1855), .Y(\myram/m6/mux_out[6] ) );
  INVX1 U1376 ( .A(n1854), .Y(\myram/m6/mux_out[5] ) );
  INVX1 U1377 ( .A(n1853), .Y(\myram/m6/mux_out[4] ) );
  INVX1 U1378 ( .A(n1852), .Y(\myram/m6/mux_out[3] ) );
  INVX1 U1379 ( .A(n1851), .Y(\myram/m6/mux_out[2] ) );
  INVX1 U1380 ( .A(n1850), .Y(\myram/m6/mux_out[1] ) );
  INVX1 U1381 ( .A(n1849), .Y(\myram/m6/mux_out[0] ) );
  INVX1 U1382 ( .A(n1898), .Y(\myram/m7/mux_out[17] ) );
  INVX1 U1383 ( .A(n1897), .Y(\myram/m7/mux_out[16] ) );
  INVX1 U1384 ( .A(n1896), .Y(\myram/m7/mux_out[15] ) );
  INVX1 U1385 ( .A(n1895), .Y(\myram/m7/mux_out[14] ) );
  INVX1 U1386 ( .A(n1894), .Y(\myram/m7/mux_out[13] ) );
  INVX1 U1387 ( .A(n1893), .Y(\myram/m7/mux_out[12] ) );
  INVX1 U1388 ( .A(n1892), .Y(\myram/m7/mux_out[11] ) );
  INVX1 U1389 ( .A(n1891), .Y(\myram/m7/mux_out[10] ) );
  INVX1 U1390 ( .A(n1890), .Y(\myram/m7/mux_out[9] ) );
  INVX1 U1391 ( .A(n1889), .Y(\myram/m7/mux_out[8] ) );
  INVX1 U1392 ( .A(n1888), .Y(\myram/m7/mux_out[7] ) );
  INVX1 U1393 ( .A(n1887), .Y(\myram/m7/mux_out[6] ) );
  INVX1 U1394 ( .A(n1886), .Y(\myram/m7/mux_out[5] ) );
  INVX1 U1395 ( .A(n1885), .Y(\myram/m7/mux_out[4] ) );
  INVX1 U1396 ( .A(n1884), .Y(\myram/m7/mux_out[3] ) );
  INVX1 U1397 ( .A(n1883), .Y(\myram/m7/mux_out[2] ) );
  INVX1 U1398 ( .A(n1882), .Y(\myram/m7/mux_out[1] ) );
  INVX1 U1399 ( .A(n1881), .Y(\myram/m7/mux_out[0] ) );
  INVX1 U1400 ( .A(n1930), .Y(\myram/m8/mux_out[17] ) );
  INVX1 U1401 ( .A(n1929), .Y(\myram/m8/mux_out[16] ) );
  INVX1 U1402 ( .A(n1928), .Y(\myram/m8/mux_out[15] ) );
  INVX1 U1403 ( .A(n1927), .Y(\myram/m8/mux_out[14] ) );
  INVX1 U1404 ( .A(n1926), .Y(\myram/m8/mux_out[13] ) );
  INVX1 U1405 ( .A(n1925), .Y(\myram/m8/mux_out[12] ) );
  INVX1 U1406 ( .A(n1924), .Y(\myram/m8/mux_out[11] ) );
  INVX1 U1407 ( .A(n1923), .Y(\myram/m8/mux_out[10] ) );
  INVX1 U1408 ( .A(n1922), .Y(\myram/m8/mux_out[9] ) );
  INVX1 U1409 ( .A(n1921), .Y(\myram/m8/mux_out[8] ) );
  INVX1 U1410 ( .A(n1920), .Y(\myram/m8/mux_out[7] ) );
  INVX1 U1411 ( .A(n1919), .Y(\myram/m8/mux_out[6] ) );
  INVX1 U1412 ( .A(n1918), .Y(\myram/m8/mux_out[5] ) );
  INVX1 U1413 ( .A(n1917), .Y(\myram/m8/mux_out[4] ) );
  INVX1 U1414 ( .A(n1916), .Y(\myram/m8/mux_out[3] ) );
  INVX1 U1415 ( .A(n1915), .Y(\myram/m8/mux_out[2] ) );
  INVX1 U1416 ( .A(n1914), .Y(\myram/m8/mux_out[1] ) );
  INVX1 U1417 ( .A(n1913), .Y(\myram/m8/mux_out[0] ) );
  INVX1 U1418 ( .A(n1962), .Y(\myram/m9/mux_out[17] ) );
  INVX1 U1419 ( .A(n1961), .Y(\myram/m9/mux_out[16] ) );
  INVX1 U1420 ( .A(n1960), .Y(\myram/m9/mux_out[15] ) );
  INVX1 U1421 ( .A(n1959), .Y(\myram/m9/mux_out[14] ) );
  INVX1 U1422 ( .A(n1958), .Y(\myram/m9/mux_out[13] ) );
  INVX1 U1423 ( .A(n1957), .Y(\myram/m9/mux_out[12] ) );
  INVX1 U1424 ( .A(n1956), .Y(\myram/m9/mux_out[11] ) );
  INVX1 U1425 ( .A(n1955), .Y(\myram/m9/mux_out[10] ) );
  INVX1 U1426 ( .A(n1954), .Y(\myram/m9/mux_out[9] ) );
  INVX1 U1427 ( .A(n1953), .Y(\myram/m9/mux_out[8] ) );
  INVX1 U1428 ( .A(n1952), .Y(\myram/m9/mux_out[7] ) );
  INVX1 U1429 ( .A(n1951), .Y(\myram/m9/mux_out[6] ) );
  INVX1 U1430 ( .A(n1950), .Y(\myram/m9/mux_out[5] ) );
  INVX1 U1431 ( .A(n1949), .Y(\myram/m9/mux_out[4] ) );
  INVX1 U1432 ( .A(n1948), .Y(\myram/m9/mux_out[3] ) );
  INVX1 U1433 ( .A(n1947), .Y(\myram/m9/mux_out[2] ) );
  INVX1 U1434 ( .A(n1946), .Y(\myram/m9/mux_out[1] ) );
  INVX1 U1435 ( .A(n1945), .Y(\myram/m9/mux_out[0] ) );
  INVX1 U1436 ( .A(n1994), .Y(\myram/m10/mux_out[17] ) );
  INVX1 U1437 ( .A(n1993), .Y(\myram/m10/mux_out[16] ) );
  INVX1 U1438 ( .A(n1992), .Y(\myram/m10/mux_out[15] ) );
  INVX1 U1439 ( .A(n1991), .Y(\myram/m10/mux_out[14] ) );
  INVX1 U1440 ( .A(n1990), .Y(\myram/m10/mux_out[13] ) );
  INVX1 U1441 ( .A(n1989), .Y(\myram/m10/mux_out[12] ) );
  INVX1 U1442 ( .A(n1988), .Y(\myram/m10/mux_out[11] ) );
  INVX1 U1443 ( .A(n1987), .Y(\myram/m10/mux_out[10] ) );
  INVX1 U1444 ( .A(n1986), .Y(\myram/m10/mux_out[9] ) );
  INVX1 U1445 ( .A(n1985), .Y(\myram/m10/mux_out[8] ) );
  INVX1 U1446 ( .A(n1984), .Y(\myram/m10/mux_out[7] ) );
  INVX1 U1447 ( .A(n1983), .Y(\myram/m10/mux_out[6] ) );
  INVX1 U1448 ( .A(n1982), .Y(\myram/m10/mux_out[5] ) );
  INVX1 U1449 ( .A(n1981), .Y(\myram/m10/mux_out[4] ) );
  INVX1 U1450 ( .A(n1980), .Y(\myram/m10/mux_out[3] ) );
  INVX1 U1451 ( .A(n1979), .Y(\myram/m10/mux_out[2] ) );
  INVX1 U1452 ( .A(n1978), .Y(\myram/m10/mux_out[1] ) );
  INVX1 U1453 ( .A(n1977), .Y(\myram/m10/mux_out[0] ) );
  INVX1 U1454 ( .A(n2026), .Y(\myram/m11/mux_out[17] ) );
  INVX1 U1455 ( .A(n2025), .Y(\myram/m11/mux_out[16] ) );
  INVX1 U1456 ( .A(n2024), .Y(\myram/m11/mux_out[15] ) );
  INVX1 U1457 ( .A(n2023), .Y(\myram/m11/mux_out[14] ) );
  INVX1 U1458 ( .A(n2022), .Y(\myram/m11/mux_out[13] ) );
  INVX1 U1459 ( .A(n2021), .Y(\myram/m11/mux_out[12] ) );
  INVX1 U1460 ( .A(n2020), .Y(\myram/m11/mux_out[11] ) );
  INVX1 U1461 ( .A(n2019), .Y(\myram/m11/mux_out[10] ) );
  INVX1 U1462 ( .A(n2018), .Y(\myram/m11/mux_out[9] ) );
  INVX1 U1463 ( .A(n2017), .Y(\myram/m11/mux_out[8] ) );
  INVX1 U1464 ( .A(n2016), .Y(\myram/m11/mux_out[7] ) );
  INVX1 U1465 ( .A(n2015), .Y(\myram/m11/mux_out[6] ) );
  INVX1 U1466 ( .A(n2014), .Y(\myram/m11/mux_out[5] ) );
  INVX1 U1467 ( .A(n2013), .Y(\myram/m11/mux_out[4] ) );
  INVX1 U1468 ( .A(n2012), .Y(\myram/m11/mux_out[3] ) );
  INVX1 U1469 ( .A(n2011), .Y(\myram/m11/mux_out[2] ) );
  INVX1 U1470 ( .A(n2010), .Y(\myram/m11/mux_out[1] ) );
  INVX1 U1471 ( .A(n2009), .Y(\myram/m11/mux_out[0] ) );
  INVX1 U1472 ( .A(n2058), .Y(\myram/m12/mux_out[17] ) );
  INVX1 U1473 ( .A(n2057), .Y(\myram/m12/mux_out[16] ) );
  INVX1 U1474 ( .A(n2056), .Y(\myram/m12/mux_out[15] ) );
  INVX1 U1475 ( .A(n2055), .Y(\myram/m12/mux_out[14] ) );
  INVX1 U1476 ( .A(n2054), .Y(\myram/m12/mux_out[13] ) );
  INVX1 U1477 ( .A(n2053), .Y(\myram/m12/mux_out[12] ) );
  INVX1 U1478 ( .A(n2052), .Y(\myram/m12/mux_out[11] ) );
  INVX1 U1479 ( .A(n2051), .Y(\myram/m12/mux_out[10] ) );
  INVX1 U1480 ( .A(n2050), .Y(\myram/m12/mux_out[9] ) );
  INVX1 U1481 ( .A(n2049), .Y(\myram/m12/mux_out[8] ) );
  INVX1 U1482 ( .A(n2048), .Y(\myram/m12/mux_out[7] ) );
  INVX1 U1483 ( .A(n2047), .Y(\myram/m12/mux_out[6] ) );
  INVX1 U1484 ( .A(n2046), .Y(\myram/m12/mux_out[5] ) );
  INVX1 U1485 ( .A(n2045), .Y(\myram/m12/mux_out[4] ) );
  INVX1 U1486 ( .A(n2044), .Y(\myram/m12/mux_out[3] ) );
  INVX1 U1487 ( .A(n2043), .Y(\myram/m12/mux_out[2] ) );
  INVX1 U1488 ( .A(n2042), .Y(\myram/m12/mux_out[1] ) );
  INVX1 U1489 ( .A(n2041), .Y(\myram/m12/mux_out[0] ) );
  INVX1 U1490 ( .A(n2090), .Y(\myram/m13/mux_out[17] ) );
  INVX1 U1491 ( .A(n2089), .Y(\myram/m13/mux_out[16] ) );
  INVX1 U1492 ( .A(n2088), .Y(\myram/m13/mux_out[15] ) );
  INVX1 U1493 ( .A(n2087), .Y(\myram/m13/mux_out[14] ) );
  INVX1 U1494 ( .A(n2086), .Y(\myram/m13/mux_out[13] ) );
  INVX1 U1495 ( .A(n2085), .Y(\myram/m13/mux_out[12] ) );
  INVX1 U1496 ( .A(n2084), .Y(\myram/m13/mux_out[11] ) );
  INVX1 U1497 ( .A(n2083), .Y(\myram/m13/mux_out[10] ) );
  INVX1 U1498 ( .A(n2082), .Y(\myram/m13/mux_out[9] ) );
  INVX1 U1499 ( .A(n2081), .Y(\myram/m13/mux_out[8] ) );
  INVX1 U1500 ( .A(n2080), .Y(\myram/m13/mux_out[7] ) );
  INVX1 U1501 ( .A(n2079), .Y(\myram/m13/mux_out[6] ) );
  INVX1 U1502 ( .A(n2078), .Y(\myram/m13/mux_out[5] ) );
  INVX1 U1503 ( .A(n2077), .Y(\myram/m13/mux_out[4] ) );
  INVX1 U1504 ( .A(n2076), .Y(\myram/m13/mux_out[3] ) );
  INVX1 U1505 ( .A(n2075), .Y(\myram/m13/mux_out[2] ) );
  INVX1 U1506 ( .A(n2074), .Y(\myram/m13/mux_out[1] ) );
  INVX1 U1507 ( .A(n2073), .Y(\myram/m13/mux_out[0] ) );
  INVX1 U1508 ( .A(n2122), .Y(\myram/m14/mux_out[17] ) );
  INVX1 U1509 ( .A(n2121), .Y(\myram/m14/mux_out[16] ) );
  INVX1 U1510 ( .A(n2120), .Y(\myram/m14/mux_out[15] ) );
  INVX1 U1511 ( .A(n2119), .Y(\myram/m14/mux_out[14] ) );
  INVX1 U1512 ( .A(n2118), .Y(\myram/m14/mux_out[13] ) );
  INVX1 U1513 ( .A(n2117), .Y(\myram/m14/mux_out[12] ) );
  INVX1 U1514 ( .A(n2116), .Y(\myram/m14/mux_out[11] ) );
  INVX1 U1515 ( .A(n2115), .Y(\myram/m14/mux_out[10] ) );
  INVX1 U1516 ( .A(n2114), .Y(\myram/m14/mux_out[9] ) );
  INVX1 U1517 ( .A(n2113), .Y(\myram/m14/mux_out[8] ) );
  INVX1 U1518 ( .A(n2112), .Y(\myram/m14/mux_out[7] ) );
  INVX1 U1519 ( .A(n2111), .Y(\myram/m14/mux_out[6] ) );
  INVX1 U1520 ( .A(n2110), .Y(\myram/m14/mux_out[5] ) );
  INVX1 U1521 ( .A(n2109), .Y(\myram/m14/mux_out[4] ) );
  INVX1 U1522 ( .A(n2108), .Y(\myram/m14/mux_out[3] ) );
  INVX1 U1523 ( .A(n2107), .Y(\myram/m14/mux_out[2] ) );
  INVX1 U1524 ( .A(n2106), .Y(\myram/m14/mux_out[1] ) );
  INVX1 U1525 ( .A(n2105), .Y(\myram/m14/mux_out[0] ) );
  INVX1 U1526 ( .A(n2154), .Y(\myram/m15/mux_out[17] ) );
  INVX1 U1527 ( .A(n2153), .Y(\myram/m15/mux_out[16] ) );
  INVX1 U1528 ( .A(n2152), .Y(\myram/m15/mux_out[15] ) );
  INVX1 U1529 ( .A(n2151), .Y(\myram/m15/mux_out[14] ) );
  INVX1 U1530 ( .A(n2150), .Y(\myram/m15/mux_out[13] ) );
  INVX1 U1531 ( .A(n2149), .Y(\myram/m15/mux_out[12] ) );
  INVX1 U1532 ( .A(n2148), .Y(\myram/m15/mux_out[11] ) );
  INVX1 U1533 ( .A(n2147), .Y(\myram/m15/mux_out[10] ) );
  INVX1 U1534 ( .A(n2146), .Y(\myram/m15/mux_out[9] ) );
  INVX1 U1535 ( .A(n2145), .Y(\myram/m15/mux_out[8] ) );
  INVX1 U1536 ( .A(n2144), .Y(\myram/m15/mux_out[7] ) );
  INVX1 U1537 ( .A(n2143), .Y(\myram/m15/mux_out[6] ) );
  INVX1 U1538 ( .A(n2142), .Y(\myram/m15/mux_out[5] ) );
  INVX1 U1539 ( .A(n2141), .Y(\myram/m15/mux_out[4] ) );
  INVX1 U1540 ( .A(n2140), .Y(\myram/m15/mux_out[3] ) );
  INVX1 U1541 ( .A(n2139), .Y(\myram/m15/mux_out[2] ) );
  INVX1 U1542 ( .A(n2138), .Y(\myram/m15/mux_out[1] ) );
  INVX1 U1543 ( .A(n2137), .Y(\myram/m15/mux_out[0] ) );
  INVX1 U1544 ( .A(n1657), .Y(\myram/m0/mux_out[0] ) );
  INVX1 U1545 ( .A(n1658), .Y(\myram/m0/mux_out[1] ) );
  INVX1 U1546 ( .A(n1659), .Y(\myram/m0/mux_out[2] ) );
  INVX1 U1547 ( .A(n1660), .Y(\myram/m0/mux_out[3] ) );
  INVX1 U1548 ( .A(n1661), .Y(\myram/m0/mux_out[4] ) );
  INVX1 U1549 ( .A(n1662), .Y(\myram/m0/mux_out[5] ) );
  INVX1 U1550 ( .A(n1663), .Y(\myram/m0/mux_out[6] ) );
  INVX1 U1551 ( .A(n1664), .Y(\myram/m0/mux_out[7] ) );
  INVX1 U1552 ( .A(n1665), .Y(\myram/m0/mux_out[8] ) );
  INVX1 U1553 ( .A(n1666), .Y(\myram/m0/mux_out[9] ) );
  INVX1 U1554 ( .A(n1667), .Y(\myram/m0/mux_out[10] ) );
  INVX1 U1555 ( .A(n1668), .Y(\myram/m0/mux_out[11] ) );
  INVX1 U1556 ( .A(n1669), .Y(\myram/m0/mux_out[12] ) );
  INVX1 U1557 ( .A(n1670), .Y(\myram/m0/mux_out[13] ) );
  INVX1 U1558 ( .A(n1671), .Y(\myram/m0/mux_out[14] ) );
  INVX1 U1559 ( .A(n1672), .Y(\myram/m0/mux_out[15] ) );
  INVX1 U1560 ( .A(n1673), .Y(\myram/m0/mux_out[16] ) );
  INVX1 U1561 ( .A(n1674), .Y(\myram/m0/mux_out[17] ) );
  INVX1 U1562 ( .A(b[3]), .Y(n1561) );
  INVX1 U1563 ( .A(b[3]), .Y(n1563) );
  INVX1 U1564 ( .A(b[3]), .Y(n1565) );
  INVX1 U1565 ( .A(b[3]), .Y(n1567) );
  INVX1 U1566 ( .A(b[3]), .Y(n1569) );
  INVX1 U1567 ( .A(b[3]), .Y(n1574) );
  INVX1 U1568 ( .A(b[3]), .Y(n1578) );
  INVX1 U1569 ( .A(b[3]), .Y(n1580) );
  INVX1 U1570 ( .A(b[3]), .Y(n1582) );
  INVX1 U1571 ( .A(b[3]), .Y(n1320) );
  INVX1 U1572 ( .A(b[3]), .Y(n1322) );
  INVX1 U1573 ( .A(b[3]), .Y(n1324) );
  INVX1 U1574 ( .A(b[3]), .Y(n1326) );
  INVX1 U1575 ( .A(b[3]), .Y(n1328) );
  INVX1 U1576 ( .A(b[3]), .Y(n1330) );
  INVX1 U1577 ( .A(b[3]), .Y(n1332) );
  INVX1 U1578 ( .A(b[3]), .Y(n1334) );
  INVX1 U1579 ( .A(b[3]), .Y(n1336) );
  INVX1 U1580 ( .A(b[3]), .Y(n1338) );
  INVX1 U1581 ( .A(b[3]), .Y(n1340) );
  INVX1 U1582 ( .A(b[3]), .Y(n1342) );
  INVX1 U1583 ( .A(b[3]), .Y(n1344) );
  INVX1 U1584 ( .A(b[3]), .Y(n1346) );
  INVX1 U1585 ( .A(b[3]), .Y(n1348) );
  INVX1 U1586 ( .A(b[3]), .Y(n1350) );
  INVX1 U1587 ( .A(b[4]), .Y(n1352) );
  INVX1 U1588 ( .A(b[4]), .Y(n1354) );
  INVX1 U1589 ( .A(b[4]), .Y(n1356) );
  INVX1 U1590 ( .A(b[4]), .Y(n1358) );
  INVX1 U1591 ( .A(b[4]), .Y(n1360) );
  INVX1 U1592 ( .A(b[4]), .Y(n1362) );
  INVX1 U1593 ( .A(b[4]), .Y(n1364) );
  INVX1 U1594 ( .A(b[4]), .Y(n1366) );
  INVX1 U1595 ( .A(b[4]), .Y(n1368) );
  INVX1 U1596 ( .A(b[4]), .Y(n1372) );
  INVX1 U1597 ( .A(b[4]), .Y(n1374) );
  INVX1 U1598 ( .A(b[4]), .Y(n1376) );
  INVX1 U1599 ( .A(b[4]), .Y(n1378) );
  INVX1 U1600 ( .A(b[4]), .Y(n1380) );
  INVX1 U1601 ( .A(b[4]), .Y(n1382) );
  INVX1 U1602 ( .A(b[4]), .Y(n1634) );
  INVX1 U1603 ( .A(b[4]), .Y(n1636) );
  INVX1 U1604 ( .A(b[4]), .Y(n1638) );
  INVX1 U1605 ( .A(b[4]), .Y(n1640) );
  INVX1 U1606 ( .A(b[4]), .Y(n1642) );
  INVX1 U1607 ( .A(b[4]), .Y(n1647) );
  INVX1 U1608 ( .A(b[4]), .Y(n1650) );
  AND2X1 U1609 ( .A(n129), .B(a[0]), .Y(\myalu/sand[0] ) );
  AND2X1 U1610 ( .A(n62), .B(a[1]), .Y(\myalu/sand[1] ) );
  AND2X1 U1611 ( .A(n25), .B(a[2]), .Y(\myalu/sand[2] ) );
  AND2X1 U1612 ( .A(b[3]), .B(a[3]), .Y(\myalu/sand[3] ) );
  AND2X1 U1613 ( .A(b[4]), .B(a[4]), .Y(\myalu/sand[4] ) );
  OR2X1 U1614 ( .A(a[23]), .B(a[22]), .Y(n12) );
  OR2X1 U1615 ( .A(a[9]), .B(a[8]), .Y(n21) );
  OR2X1 U1616 ( .A(a[30]), .B(a[2]), .Y(n23) );
  OR2X1 U1617 ( .A(a[16]), .B(a[15]), .Y(n14) );
  OR2X1 U1618 ( .A(a[12]), .B(a[11]), .Y(n15) );
  OR2X1 U1619 ( .A(a[27]), .B(a[26]), .Y(n24) );
  INVX1 U1620 ( .A(n1512), .Y(\myalu/mysrl/s2[31] ) );
  INVX1 U1621 ( .A(n1608), .Y(\myalu/mysrl/s4[31] ) );
  INVX1 U1622 ( .A(n1560), .Y(\myalu/mysrl/s3[31] ) );
  INVX1 U1623 ( .A(n1464), .Y(\myalu/mysrl/s1[31] ) );
  INVX1 U1624 ( .A(b[0]), .Y(n1463) );
  INVX1 U1625 ( .A(n959), .Y(\mypc/temp_pc0[7] ) );
  INVX1 U1626 ( .A(n954), .Y(\mypc/temp_pc0[2] ) );
  INVX1 U1627 ( .A(n955), .Y(\mypc/temp_pc0[3] ) );
  INVX1 U1628 ( .A(n958), .Y(\mypc/temp_pc0[6] ) );
  INVX1 U1629 ( .A(n1010), .Y(\myalu/s10[9] ) );
  AND2X1 U1630 ( .A(b[9]), .B(a[9]), .Y(\myalu/sand[9] ) );
  AND2X1 U1631 ( .A(n10), .B(n11), .Y(n9) );
  OR2X1 U1632 ( .A(a[1]), .B(a[19]), .Y(n13) );
  AND2X1 U1633 ( .A(n19), .B(n20), .Y(n18) );
  OR2X1 U1634 ( .A(a[5]), .B(a[4]), .Y(n22) );
  AND2X1 U1635 ( .A(\mypc/temp_pc1[1] ), .B(power), .Y(next_pc[1]) );
  AND2X1 U1636 ( .A(\mypc/temp_pc1[2] ), .B(power), .Y(next_pc[2]) );
  AND2X1 U1637 ( .A(\mypc/temp_pc1[3] ), .B(power), .Y(next_pc[3]) );
  AND2X1 U1638 ( .A(\mypc/temp_pc1[4] ), .B(power), .Y(next_pc[4]) );
  AND2X1 U1639 ( .A(\mypc/temp_pc1[5] ), .B(power), .Y(next_pc[5]) );
  AND2X1 U1640 ( .A(\mypc/temp_pc1[6] ), .B(power), .Y(next_pc[6]) );
  AND2X1 U1641 ( .A(\mypc/temp_pc1[7] ), .B(power), .Y(next_pc[7]) );
  AND2X1 U1642 ( .A(\mypc/temp_pc1[0] ), .B(power), .Y(next_pc[0]) );
  AND2X1 U1643 ( .A(b[26]), .B(a[26]), .Y(\myalu/sand[26] ) );
  AND2X1 U1644 ( .A(b[27]), .B(a[27]), .Y(\myalu/sand[27] ) );
  AND2X1 U1645 ( .A(b[28]), .B(a[28]), .Y(\myalu/sand[28] ) );
  AND2X1 U1646 ( .A(b[29]), .B(a[29]), .Y(\myalu/sand[29] ) );
  AND2X1 U1647 ( .A(b[30]), .B(a[30]), .Y(\myalu/sand[30] ) );
  AND2X1 U1648 ( .A(b[31]), .B(a[31]), .Y(\myalu/sand[31] ) );
  AND2X1 U1649 ( .A(b[5]), .B(a[5]), .Y(\myalu/sand[5] ) );
  AND2X1 U1650 ( .A(b[6]), .B(a[6]), .Y(\myalu/sand[6] ) );
  AND2X1 U1651 ( .A(b[7]), .B(a[7]), .Y(\myalu/sand[7] ) );
  AND2X1 U1652 ( .A(b[8]), .B(a[8]), .Y(\myalu/sand[8] ) );
  AND2X1 U1653 ( .A(b[10]), .B(a[10]), .Y(\myalu/sand[10] ) );
  AND2X1 U1654 ( .A(b[11]), .B(a[11]), .Y(\myalu/sand[11] ) );
  AND2X1 U1655 ( .A(b[12]), .B(a[12]), .Y(\myalu/sand[12] ) );
  AND2X1 U1656 ( .A(b[13]), .B(a[13]), .Y(\myalu/sand[13] ) );
  AND2X1 U1657 ( .A(b[14]), .B(a[14]), .Y(\myalu/sand[14] ) );
  AND2X1 U1658 ( .A(b[15]), .B(a[15]), .Y(\myalu/sand[15] ) );
  AND2X1 U1659 ( .A(b[16]), .B(a[16]), .Y(\myalu/sand[16] ) );
  AND2X1 U1660 ( .A(b[17]), .B(a[17]), .Y(\myalu/sand[17] ) );
  AND2X1 U1661 ( .A(b[18]), .B(a[18]), .Y(\myalu/sand[18] ) );
  AND2X1 U1662 ( .A(b[19]), .B(a[19]), .Y(\myalu/sand[19] ) );
  AND2X1 U1663 ( .A(b[20]), .B(a[20]), .Y(\myalu/sand[20] ) );
  AND2X1 U1664 ( .A(b[21]), .B(a[21]), .Y(\myalu/sand[21] ) );
  AND2X1 U1665 ( .A(b[22]), .B(a[22]), .Y(\myalu/sand[22] ) );
  AND2X1 U1666 ( .A(b[23]), .B(a[23]), .Y(\myalu/sand[23] ) );
  AND2X1 U1667 ( .A(b[24]), .B(a[24]), .Y(\myalu/sand[24] ) );
  AND2X1 U1668 ( .A(b[25]), .B(a[25]), .Y(\myalu/sand[25] ) );
  BUFX2 U1669 ( .A(stop_en), .Y(n211) );
  BUFX2 U1670 ( .A(addr_s[0]), .Y(n209) );
  BUFX2 U1671 ( .A(addr_s[1]), .Y(n210) );
  OR2X1 U1672 ( .A(addr_s[2]), .B(n841), .Y(n203) );
  OR2X1 U1673 ( .A(addr_s[2]), .B(\myram/ds/en0 ), .Y(n204) );
  INVX1 U1674 ( .A(\myram/ds/d0/en1 ), .Y(n837) );
  INVX1 U1675 ( .A(\myram/ds/d1/en1 ), .Y(n839) );
  AND2X1 U1676 ( .A(addr_s[2]), .B(\myram/ds/en1 ), .Y(\myram/ds/d1/en1 ) );
  INVX1 U1677 ( .A(pc[1]), .Y(n842) );
  INVX1 U1678 ( .A(pc[2]), .Y(n843) );
  INVX1 U1679 ( .A(pc[3]), .Y(n844) );
  INVX1 U1680 ( .A(pc[4]), .Y(n845) );
  INVX1 U1681 ( .A(pc[5]), .Y(n846) );
  INVX1 U1682 ( .A(pc[6]), .Y(n847) );
  INVX1 U1683 ( .A(pc[7]), .Y(n848) );
  INVX1 U1684 ( .A(pc[0]), .Y(\mypc/inc_pc[0] ) );
endmodule

